XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>t7s�
�7e���zӁn}^�iu�B���Q-9Qi�ܸHk�N�Z�l�$V1�|�+��A�"v���cEJ�g�g�|�O�1#^�2�E�K'�h�6<��;��Y��%ݞ�?����Q����a()~n:�K.�q�����*~�o��F�:a�Q�/Ҡ��
k����j �������<F[q��oy����d�9�`](Ҷ&cǪ�7=ԛU�����\� �Bς:�8����J�f���U�7�[�y���G4�-y+c0�'Ee(����g�/\x4�C���� \&}	�,<�h��H��
�
�>��l.R�w����� ��C���}&S�y��Źf�)ӶN������:��';��Ȥ�"�i�N��K��I�tǻU��N��z$*��}^�
y�����T�ō�Y��H�S��_XX�i����,b_O�v�B�{V�L�h�;�L/��)�N ���᥎��U������Yt���u��s�.L�:��@�����1<ќ蓕��"�{hg�3Zhl�-�!��aZ�����5^�r�$0(gF<�f�*�я�<f�{c]��6��m0���rUY�>����|��v�I,`�G�ཱྀ'��Z;j�ZT��9�l�o�*o�,W��"s��k|E�k�����$So�Dx�\�քv��WVn�;]��%���=���Kg� ���V'VE���+��8�e����?²1�e�|K4�,<��)�C��|`s��>$x���"XlxVHYEB    55a7     e50j���%�x��8g�?E���#�"�(�;�~7��$����*�#��>ȯ�����ܘ\�m���9[`�&XYIuO��,�ZpP����ԠpIH���S>� ��ˎ�C���9l�r ����;�<�K��O��b��j����oK�uj�q�B	Pb�->�����3k� ��Ä�vZFW3�����������O[А��&���u��{���0�9���x_?��b%���Eg�����k7�Pŧ��g�) Aښwzk�oR�l]���4�=Ȱp�,<�<|�c?$9P	A0S�s�\�x[����M �1VE�Ȕ���1��dw�|�u�����h�������y��;�EX�AZ����ʩ�#�9ɼ��8�?X=:�?�"Axf��+|�l�	�"Q��wغMaO�Jť��#�	U~�î6�ӄ����~�OO�0�HKx2[(o>	[��e��r�'Yeh����ko��N�"�%�!Q��WC��G�.*�ͩ����鉙�Rׁ�p�=�	�t$���~�[F<��5�C���v���k�5IV�l�Z���$"�5��x�钔v��^��tC��\�PX��ك��(Otb��,P%>��m=�i��9��{!�H�qY\��J�w��魕���N�C ���M8k����ى��&(-�"�(�s�}��hN�E��m��&(R1��G�}��3PQ�����"3�"A��墶�}V(�'9�	����k�+�ÿ�30�Ţ|}����]ge��1,�h��u�s�6�ZKpT��s�=��zQ�=^�<��Ss�R�h�	nrqnP9��CM���D��9�nF77BZ��Y/�'��ŴΥ����W=�άSz��h!3���b|����a(���:�qvM��ӵ���_�W�?.��P,�y��e�`l7"Дs�����G��y�{R�@�ԃ���X�V����n��x�d?��ȭ�U�e�G�7�-�����ՙ��v�輛����cy�Wx�:�o��礸SR�g���:�r��鱶xmO�5F�<@���X�-��o�9S�#�&�n�j���`�C��{���w����b��9A��J�ƍ�x�J	�a��*"nwA~���	�ݻyX�r��L�d�[�^Gv\��m����d��i�@�N�jgc�2�>�1)�~E����4��s����#.��ʿ�8���f$R|���p�沤�K����P�뒥#�E��=��}&FQ�R�d��|uzÚǌ=��z߅�ী�c:é�����w{(G��Gr� H���������)_|���$���W5j���T+�����~{�դ܊����M���諙[�0�̄g)�=QD�4 5-/C�"�-d�C��C�ֲ�����+ ~xzT�y�q��6,ϑ�@B��i�W�����v�>����cj�M��^�y�8V���46���TtfE��T/��20��x:��"��@�r-m|�SR�?���J=ˋ�Ra},!��3x{���q����>�o9�J�:W҄�����)Zt�DY�e��O��g|?2�M�#o�:��N�OQ���|P��a����2�T���k�\�y7���U�~&��҄"��m|�������J�=X��c�O^����@�ŷF�:j��|_N�p���QfC��2JNR��i�'3	79���qI����$���x"ko�y+��Þy���5(,�R|M��*�.ZQ�+�3���6�@Զ��m�0����H�a�\{��������+�O���pͼ�l�����D���x0�z序n!����9U򌉢��6&�c�o�m�!�|*���_�.��(�-iyI!�&go	U�d �M&ȅ������b��?)��[�+!f{���H	��wGsMj憹�?�#����X�<���c�_���)8����]�!,�\�uŶQ������'�\���H�"mb�e���1�5�=�)�p:I���4�廰T�H�},���n��џN���n�R7`B��z��`��l�[��������9嗗��=������0�b��m��x��L,�	�F��n@��
����P�6�Cy�bƜ�;�YzCb�i�z]�_����{���*~+Um��ո�r�B]��$����VQ@�g�~	��BC���9�d�T2�O����k�/�+5ߠh'��>�Jv�J�ʱ  ��λ��j�p�~�c�W�i�6�;i��lkG<6�6;�N6��:t~M��T�5͎~�Q쇬h
���&=-9�x��6�?tƵ��!�J��jr���^�C���q�Xn�ħg]�;ok_mQ��M�wʊ�k4k�xQ���1I��$~	�K��"SNAyk��5 W>^7�º2t�3��`�x.pSF�p樉�k
!'y���r �_	F�µO�1	_ހ�m�­E�~���'��'�.���*7E�6�YN\�q<f�G��A�Ϡ��h�n����i@Eؕ7G�^��Yn�=R���b�=SS^}����L+t�$8����=��]m`E���Ne�&	�ۏف�p���A��bQ�B���6�8��Hl���\tQ�2O��u~�+O�*:�2�_�1$u��vix�Z�d9$��~aTc!K�N~���{j�,���v����Vg�~ϒdd�);E.u�^.i,���*Z9�g<�i�A�Gh��a��&(E�������86ή1���X	(�W2��\y���?6�+�2&�옡4)��}k�z	���T����r�CN�R�=_�	גf��TR���L����w�4���}����ȧ�ϊ�h���硆����$����_(�˖?�8�!-�luO��_��*���2�� s��Ӊz�;��X���
u{c/05���e.[�˝�	����Ƃ��n���a߆62[~�ܹ7<R[S]�Q���|��� �gۢ�h�b#*� �(@�NfS8�a��G͚��es6�����
c��˨΅�Ϸ���!]򪣻é�����+�=�ޞ��ˤ
|0��1�~z���'-n��:W����'�v�����$��k̚34���A�"�|o��Ʈ%�m0]�W��(	sJ��h�w���ph�'�2���,���N���(��FKlH�,���8�4�ω��~�Y?��ݶd�Ԁ]�uø���R�f�����S>���"��x��wh*�����J�ኊ��qy��ޤ��S�}��=���軱NY�Ob8
z�[8�yn50�u2�qsh��#Id��-�.�����������}�A�L)�>�/�[ӝ'U�kn�݄}�3tK����`������(�i"(��e�����#O���tݏ�C���(�;c,�I3�e�j�"L=\K��� ���*2�oȋ��Jr	�a�Wf�a��&8u��-5Y�Y�OF��5���/xG�_H�fh�pm�٬�7�4ܩ��ӣG!Z��~]�K�jS�E��G��ié���%�n-Z8��SV/|���L^/���\3�Y�4>��F�&��d0�<>�U�J�����UOI*��YS��Y����M�]]y�Y޷�?�����a�hy�6,;ՙ�U�5�b^i��ȣR��E�c_s����|���