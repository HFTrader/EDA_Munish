XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��E.d�'�A`�=�t�`�X�N�����rL��=e�`�'���tr���T����qm���1�L������L=G.|�4p��M5k��,�#�3z��O?�U	}/u�v�!5ŗ�|U��9_�V~�kq����/bN�*�0��v�I�^�Y�y	�pJ?#s��A��,n��A��Q� v�W׾�E�o5P<M�PR?�RW��¿�G�������<aC+n%Р`�k�z��
�J5�����#���Q4���Bi���>s�^�iJ�7X���@=j8Ʀ9���%�v����Z:h#X��	���HX0e��MqҬg`R��0|� ���&�:�^��h-.���s�"���%���x��FVI�*�}��p#����%�<�m��k7_�ag�Ҋ�����P4��=Yu+�����ПE�$gI�� N��Ĵ<s�5t��sǦ�:/v�Ag�_S��֘O��@	d*�\<uAirYK�Brĉk=K䕍?U�<m/�k�L`��d�--�p�ի�,�\[U�?��J?*|툂��(
7�􇌌�|������
e�9zm'��ߣjkO�p�>4��0��"&��B�L�5M9W��xr+X�q��JjUtA�6���[�D�_\p:Y�k���R>0l���Qw~3�hN��}��A�7tZ�0i�yc�R�2����b��_'
��?��]�C7э�z��<��$�f�W�
'4�c▊�L�_D�Sl�\���b8 ��XlxVHYEB    aa31    1e40����*ox7���IE�y��8����
.�T[R��(����ȭ(u �EC_B���=@��S�_q����z^��s|�iZ1�$��7n�p�
�9E7q�0U�������
�$b֦Xp^�HW���d�,� 7CMD�1݉r�
=�K�W�\�ۆ������E|[���~�v��_ �����dÙ�?qc�J %�-Y��~?�E������R�3.l;��L�4O���;^�Wμ��ҏ``��5��k�j�߁������7��y\�d�x�;n�M��^���|���Μ��KW\��s���3�ͅ��K	s2��`TP�E�I���DҀa�CJ�@y1O�2�D�5K��� ����pC�h�a�ڰ�?h3�Z����6q��$ �>�~�|3���Q��.l!���|ys���P󒂧s�`|�KZ��{_�ރ:&\�ڪ2Gw�s��)h5T֍�v���ԇ׼)4N���K��_	.v���&j_A6Z�̗W����񻱠�ѺB����`�CF�4 ����t�oO	F`��TB�%ҜZ[.�	7zJ��݊��EU�4���������1&��"ߛ�.?�z0la ח�C)�2,g��1DS�"T�bw��:pA�-[b�<fߩ�um��Q@�Pl� ڞ�!�A_�n<���
맋�K���y"�u��ǫ�#��m�b�hw�iUZb�V��
�	�!�c��"�Ԥ��+�
҈�"+� G�:�'D[�eVM�FjX�����?����E��s���믮�ɲ�..�+�>�\�:D���I�:��y_�	���S4��g~���� $������{�8U����-���X�w/6$����}�]Nh�:ݲ�P.���_��ږ�n�b-Ѵ=�0+� ������U�'�~o��bY>3	�]�b��`���cx��.-=# ��^^TK��3�Hy�yjma���+�F��	&��l�,�?�����@g[�I�;��4%~㊪	�g��B���T�|�IR�д����߿�w�^�׆d�+����`s�E�O����2�8v�I�Ds�\�N(����Ε�B姠I�R\�$oIܓ�v��ʹ���n9���2K�¤1����}.l��<:�k2�'��/�jnS���oA���ꗌ͋�Ӏ�O�҅|;������-���ܣ�a���N΃"�a��ޣ�@�^������~�:�ni����N�@T�%��߳ZL΅C����~%
 �s9<9<H�}Obt����3�o��,�2�8���������,4��`�rT�������Q�L�-y3:����eN��Ր��0��50���o
��[k(f�1�t�h�z���c��lUC�!4���-�@����P�f	c[$6X=/{� �?��t��o��h`-�Al}П��&�-'�z�Fh�҈΍zR���tY%�5�Ye�ٖ Y�%�<�-4��:\Q��)C��*���`Sdװ㸃R���5B%�eC�G{]��ܙP�2��p�T���ފ#��{�x��C�(��PCnN�G�gqɸ�i|x@ �.�F�E�� ��-������v��-�t-�ȫ�ܚQ]8&�Y�VmdF���bO8��F<I���5n��RB�����uX5jE٭�su9b^�9ҡvLg�����H:�,��n���wv!8	�A[���>���q��a���'R(bhʾ��0)��KQNup���I��K;D�3I�\�L��F3���d�UЕ'���8�qb⃄�D�R�}{�ѾE�R�ob��^�,/�Mq��VŐ7���M#úU�%a�5-Zw>	w�/��?L�,BoJƻ��Ԟr��[�I�7K�K�̯a���J�l�_T� 8
?ۑ�F��vZ���0��N
D��ZW�룄��	�ۉ-{#U~�s��#�l�*\瞗L(5R����;<ߥ�p>-D= h]C��HE�\A^h��.�י'�u���}����<�f���C/%���p�Kr�������.�=J�������I�q �,��@hr>^V�6�R�~gi��wĚ<Q'�yy���)Y>����ԅê��M�z��R6ꍁ�p�H�bl�D+�i��y��4��<׎���-�U��}�h� F��9� WԴE���Y�W��#���7�q��?h�u����'�<�AR�tG৤y�ϱ��D�����43r�,��]�"(	���~������Q��u5i�'<��'w��&�?S��@��	�$�� ׎A���|������/n�T�=�-�8y���=���[�k��^����M�+E�RwLH�� �!k�[:��~��\*����H4bզ��04��ۓ�]:-��&~�O���7��0e�	�蠻&E���)�71K_xk�iS�*ǻ�[Q�.fQ�����7l&4b7��N� ��>a�����$!~�a�4~h�h��dn��ud��,���3���"�t���O<���|�
�偩v�����2�7 �F���F?�ˏJ!G%�u��9P�J�=C��;��������Y��O,������X7�%�A�#x\ֳE g�0^R�����U�Ά�O�������b�����̀f!�-�6g�%1�_�A��'���~�"��2��'����p�/;}��:�Dп*���oP+3+O=��}��e�;�=}�(�k��ݾ���H�$=C����Tь�M�{�1R-�	�6�mTZ�l�3�S��|ܾB�I{�����Rt𶂔�&@@�=�/�T�"ũb����gnt�x��%��Ðzݑ&椏�/��˛3��c���mܰ�,N��F�7
�ֶ݉��2>"ֽfc�9!#�3�:�<�������3j�A�	eD�&�\.�l��<p���v�L'|�g�9UЪ���w��ol��|_��KM����哌ܽ�B3�k~UddG��9���3%g��;���*-Ǽ^ͼ�pҰ�����~mHl���uѭKk�A~���E1&�,w�v�O�|@��t6_9��rx�z�E��\�?X��֟zB�C����%%�]a,-?|V|&o�*�Yi����mo�ɀcy�:l��߄��3�Eh�}C��	-s^�͆�����5Kk�6�"4�nC�/2�}#G�~��U,{dA[/n-Z�8x�h���� ��������pT���J%y9�^S��Ϝ�S~�K��W�79Wnha� �U�����.E����`��"1%iu���V@�� ��)��ӛp��y�4Ԏg��U��M�CHf�52i};[$\�!�!��0|��M�՝�/{zG#td_�cX�r4Π���T���A�b
͙-2�_:lZ�փ�:��J���C�O���ql?uт-�g�,U����.��;�|a�`/�`�>�:�O���\w��DP�=pb;l4p��6�!�2�DMAt1�dCbX]���-��Ʒ���K��ijc������&�*Stdc���Cş�?���Nڑ��ۼa�0H�鈕,	Rs }�ـW��w�r�9����Y������

|��DL��p)ωB�ON�@�M��J�a�9ı��U�9	6R4�g�q��(:7����uҺ�@`�Њ�z��ۺ�ʵ�3�z�s	���:Ȭ�m}���؃^f/J�����ksSn�4�W���c#�@UO��kE0�Ab\��P�;t�2�I����<�"<L�x�Nh��AF_�R�����7C|� ��Lȟ���5C��Nly!����e:�j�u���v��y�?����J���L� ��~i'ƣ�*���As�Hag��R�0	��� 4r)�i���飶�������� ��p#(��t�L��ӯ7c�p��)/zu�f�"�6+�����7�
�c�N?8@E�R�"���S\ o��(r�Kz�d'B�sP��¾��z:I�jt�1}r=�(�,M4���}]J�Iz�&��Z;AZ���ωy���M��y�x��I�<F|e'���\mm��;��sy���S��K�=��O�����^��	l��,�L��GnrN�K�>�1/���&	�r9��C�8w�N3��p���ƚ;�x���P�Lo�v@8��M44q�RF���X�b>�@����3]b?�8@�8�n�����U�˒Nȴa�*(�RF_�Je�5L�E��J�y����W�g�!��d�?�-�9��|��g4��"g��?;��iv4�N9�8�|4�~�Z54�'6��OI1\=��B�d���9v�z�D_�����޸�SK8¨䷠��F�����||a'��?G�}����a�]�\�u���G�)���:��%s����O%z8$*��+FaX�鮇E��M?�N��.ڹ�%�~B<�D>�/\��m߮ �ɵ�y�c��H\��{/�Q����~CȏΕ��x���R�ԡ����h�Lȶ}��n�ZBW���\���� �$�M��]�=ᄺ�R���лg�uf�DN�p[�L]�Bh���2�_������g��nOUx4�h����)��Y�9��4���b0�c��׈��"��i��2{8������'G���A�Ҿ�ڜM�����c�)_e���W�|���p�I�۵x��,#�佻���`���I�x���\��(����j�Զ1��"2ܿO�~M���`^��=,y^I���]�1pmU��Nߍ���2]�u~�m%�����:�}���k�/�����6VH�f��n�fB��O���<��EAyz	���kˣC�F�&��v��Y~AV,�6a%��OCl#��������ـQYW�>MY����G�v,�	�~�D���k�[��}�*:Z*��+�ާ����N�Fxi�b�x��m���OU�	�H}��c��݋oO���6rJ�OS)�M���N�����tH���m�ȡ^�T5ݠܑr�c�A$0s"tw��6�٧� ��Š>5*:?��/���&?�������~���`k����ٝ�f`߻n���� c�(��ٸ�V:�;k4��[��p��3�k�����_�C��F8~({E�^�#�9{<���vz3�g�-�~Ȧ���&d��(w3��Q���勃�n.�BvM��\�+��>fʝC
�!8	�rQN�[�<��X�Ĳi�)�Q�����T�l|�p���i~y�7`�V��~7pB �CT۸�L��8���e=�<f{���P�?�3V�~r1��uv;W��V��9G��GM��u2�<�=j>`�{�EPu���}�R�c[�CH����[ӚJ��������T��E�x���{��%��R�?�q�`UrAś��Lm���# ��C�V�4�>g{�'��G��{��d6���ӝ�*�髆��u�oR�
��i��K���OO��/"A3~z��H� `J��JV��W�qCC�y�\�3tG�a�{>��Qǟg,.�]�_��gt&�Vq��ϑ�l�#!a�s>��t�HK	 ����D�RQ�,Ǔzǁ+��R�}|B�g��m���~J�b�_y�ZL�����&/�H����n���L���`�������R�Ob�&��Er/y����1������s4��;�{�?ͮ���z���Q�W.���:�!�-ќ�s��՟�_	�6�����vP oo�pM����9�w��mek~�ڂ�t���H l{�"��Vi`?/:�j�V�����D��.[����S������[���܉]y���fѕ[dg[A�F�`oI�I����n�NI���`s.��4������dz�d��_�����r�1�9�I���V���;H��� ŔA���2u�B����TąD�ik�+��5+r�GYX��,�qp��FM�Hç)�ݯ��#Q�;�TyZ5$��m��X�1�!�TbQ����(�f�?!M��EK���S����w���jP�mbYf��;�sQ��k�L�Ltw�$�<�_��8Z�q��ߠ�����XT�{�fÉٓЀw�'�uY��e���m8��}�����b!�=D�<���1����K}�Bz�i9=Q=�T�Z�'�*�؏�y+�I%]�2�ky�l��6�K�(���$�J��#<8�q�ч��!��AX'0)�铌��ũ��y5#��ڻ=}^�U"�:��>� �p� Q`r>����_��#���9͑��șjF�=�r�k{��l�s�Gv8�4�GZ����`q��Dc��r�!��1`���$��:�Yn��:����+���N������p�
܇�lYH���þ���8޹�R
���ň=EWD�O��/6?�]T<�K�qՙ�D�wV��Mg�W�3{C)}o���/�7u(��S���;N�[uR4�}���Q_�m�M��&G'��Z|��V�|��oMI�'���e|l�8J��K�17eq��F�]�[&d]��{��6~R��Eɪ��}��_�`4KJ^�u�vi��;`�>@p�(q7G�4�Rn��g)wa?��ĺ�z�eSVޫa@���@A�&{*%�(��XM1��->c(�Xع|�	^����4y��>����;�!�.�3+��^?�ڇ��xK%T��V[�'��I��d�x�Q�,��#L�gZFWMd�^v��\�m�X�e�o�X"(�OFp��f0B);��m$r3�Ĳ{J�ryH/�����M �H�VΨ���(<"���|�>U.�6�w^$+�OC�u�ӏ��m0�ĕ�3"���_��˥�w�G0Q��oYq�>�.��Ԑޱ  �N�(���X�de��Оl��gA!��\	
w�T#��sz��K�n�����h^D|�!��LF2} �e�h3,`�</O�·^ͻ�1������y��#(�"�q�u���^h���P�^}�.������#�A ���~H𙟉�L(dl��5�l�{o��m0�p���(�]۵Ч�ٲ���Rfs�� �O�8��0x� ^'p��~������DeO�~�PЗB�Kp����;>
�͒�.�~C1� Vm��_@a��Om�?��e�EC�m�������ED䪏bU���NJ~�x�)��:�Ň3�}z�o]�7�̴���ϴiݮp�* O,P���G��&��:T�+�?ի^,��B ��B=�(��i��!ּ��yg �
Z�};���$�����?��tA+B�e�
S�/�:���P�o���^�l�E�c������Gm.!�G�@?��a���T�v^f��et�_yA3X����P}S�Ehе����"+설�('1 J�<߸o fY��v��X4��wg���.���|S�I�|vSva��{[?��)�X�s��%J��d�Q�_���k���m$��H{������`�1e��=������|�_�]�L�n�	6_@6�IF"*	�Cui[��aHB\J�A'��8�to릓��3�N�.�p���{�3Xc��.����H</Z�q9���I�
���*ST���V�<�U_�zO���`T.Z�M�R�=�粎� �]�0�S�A�YR
�ą���V��: I����<t=�!����S���T�p��
>; �N��R[=!�J����"�(}dH����m�?pR��m���S8u'^Y�sEA��Gc�}~