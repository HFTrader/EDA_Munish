XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���*�9p�:�.�[� �����P�*���r��.j�HBs���\��p�R�����,q:���O�݈㤤}I�Γ�;�r%
�E��\�]FC��� t�vv%m�%��,��'�ί@�d�
eT�c�2�ܪ��P��"HxŬ�Z���n�l��O<"<�Bk�u��BF���z)I���^8�X�Ux�oE7������/�-�/��x�Ct�~�5@*��ȶ�_>��@[v���;q<@ϳx�}��g/v�T➰�\G�����Q	)YZW'�U�`���9䉂��l|z�c�P�j�سg؜��e����Pe���,	�P�bL<���0\ᅒ�@@!���o��� #䝫�����I�z_6��]08H��a愡�����Z��(��������C��
)�����Q0�Q{�L�]ܺ�����9X�hݱ���1A��",�C#*��?�s��2���ɺ@��#~<�������3�k�9-f����g��G@v/�=��Js(
<��uV.y�ի��������o�OX�u~m�~��i���H07hm����in+ԭ�y�J��G>�C쫪ï�����>���E���#k�d�F:�@�iй����j�slF*��=m[?CnW�x��-&w�����	����>£a�o9�nɱP��mJ6̽��� 
�GƋ�8O�6 V�==��K4awT�x�U��>,.�������0��nv��ԑpf._���P�LQ@�U���nN�a�c�A��XlxVHYEB    fa00    2030g�w�Վ���^��P�#��B�ԇh���3%z#�P ��� �pڠ[R�'�^;�,�����M�����n�����+�G�_�zO�>��"6󓖆������uS��@�	������jx-��
�-���_7$��> w��g� AFHb�*�=}�Q`��~��1y
��o?��+��|E�A$�\�����崥��`��E�=B��!T,.� �f���<O�>
��<X�Ġ�	���g������V��f����s��I��z] P؅���t�Dt=�H�Y��wUÌ@�Kn�u�ҵǵ1���3�!�Կ2�_2�ш�`S��[DEyuj%]��:�ј1o7����8�/x���)�����D��������F�g=�DQ�������A�����%֕���^8s�U��su����G��J���\�[I.eV]q@8��x�-��.y��D_�����ϡ/�X��vSx9h8=m��X�
"ͪƚ���s�{�]IZ/�����y�/�W�l*��!� ���YF����f��X�X<�8:�߁#������ǻ<�K� �]�����E*��8n$����_�i�#w�D�In�t!G!%��5�r���C>��M���HdB��Ġ���z*<�Q#���P<yg�l�ݿ��K�EÞ'�w�Z�����k����?����T��$��N�o��Jz�l���3ƲUb@f>��n�J�+���e�_m�N���r�)Ǐ#_��(ܭ��o7�5sO�/8#����?k�X>����ci�k/���=_��Um�!.w��ЖP�Nُ����aG�Nq��oL��x�C�^xuV`�~��_�Q���*6�eTp$��]�v/YU�--�k�f��*��W')��㨹S@1��3Q��\��iA����4Q��e�@�D(cպ-Z� ��o˿�V�R����L���pRt�<?DQa�ὲ*L������@,�h8��)<���ݡ��4����T�20jÿ���ۺ`:��0��=���m�B>��7��=<��>Pԛ*/�2�"Q=YK�Cq�՞m�G�_�:2|^��w!�)(X`���Uft�)�su�7��Y��v�=��l�"��>�:���U>�&���߯�o�d[4��d���_�Qm�	ET���`��:�9��&�z��u�@����T'�����p�hJh�j�n�>��]�4�=+e!@Qц޺5y%pOY�=�4[K��:��?N
�Bi����S��P*�F!�YQX�aF�:�JrN��.ָ~�o���������!��V;?�n��l�@7�A('�u��W�J�;�gjO�IC�%L�DO�KZ�:O�yͬ�賘 ���u�lF��ZȨ�IGЗ���\a$���C.jtv*_!�:s��v<�\��TP"5��/C2��0/&������Ӷ���N>�R��m�k�/p���BP�Dx
;��CdH�+�Ӈ.K�+�Q��?B̂�u��4�u3����	����2=��@j���ћ������.��s-gE:�F[�i
h[����:<���$L�ǀ� �̾�^��,ZrLs��'�����T���Čjt��tAM�)B���ϟ#UN�	�?�n����rNp�:�6�����ymְus(��y0�%%�(\du���a����@4�.
���:c��:Y��m��t��ۀpy�)9��4�шb�LX6��"��(��TRc	�? ���gg��E~?��a��7�'Qϐ_ݯ�2gV���e�������a��\�b+~�~O�|p����H��ߔ,\�h�ı��`�4������ N	��d�9�Ow�Tj��x�E����$�������x�T�]O��p$��g��OZ\i�"�H]���]�[H$�L�����J��6��UN�B�����d��I�v`?�ϊ� M4�I|r-�����J��#v���hZjZ*�5!��G�/������)�y�h� [5p��E�E�Hܙ�\䒝��3���5���Ϲ��!�Ҥ/Y��]���Ո6=]r��5��*X
�~���Ŧ�L��q�`c+6x��fIE.��:l��+'_�<0s���l9�#7A���o�R��p���//��ks�i9WЖ6 ���[4�bONL��?L�'��2�K$!�<Y��=�������\��U��-#�Cw3���F��J��sN��$�0E�#��l[x�-��������eI�f�߉qAl�`��6$��W�h���\&(VW(ۣ:�\g2��P�v�����(Խ�F�Q���0���_����{�%��/�y��e�;/��4W_�oG��+nĹ��g�պ!�֥��D��+�φ�h��A�2�`
*�1e]�>.}�� -d*�\��>��/+}ʡ�����7i@�'BU1�\I+�@X�}�M������_>�G���xw�⳨�>2�w7Wذ�����#ѴRs����v:B�SD��'僓�VMt�Cޢ�8B�pf���0g���K�x�A��L��%��֗��7?�*�AKkP�x� ]�e�X�0=�첥X��Qd�Ԏm9;y068��p��A.�^\� �zo�<�o��^�3 ��U���z��:��5Ф�4mtc�Z��I�dNA�dr-[��.�ϯ�w�w)o��e���o�[.�>���#e�I�q�h&��G�K��C��N>���q5"p����|��f���ϰi�R}�{s��W�[W�ӿ�P����w!����{�?9M+|_�}���T���Q�D��_���@��|t,��pIT�_�� Ӈ�o���F�S��-?=)Õk�i�G�Sg����������NY	��0��yX��;��� �M8תdp	��_�^���)���6�6 |�8HO�o?��lǠ�H��H���e�}9Lc���틢��e�&r2��z��d��[�h�a��+�؁n;����(�G�/'+[k�[��99S�Ã�#��q��ӶS�!��F��d2Ѐ��S3�5nJ4���"U�[��1��S�30i������4oVC$�o��g�����V�P�g�w|8�9ٞ�V�[JV�(s��c>�lƘ���M�Y-xۘJ��/u��j:CD� ���j���x��I Ld�$n�����N���E �r${L$#�NQfj���cˌ#�@P`��T�4�:2s2�:� ���D���d��&+DLg.��m��#�Z��<��aY��V#��#��� 6���=^�#�zR�&���ƭ�,���O��[��P �l�wi�w�:2���8\~	as^��c&3d�����n@�m����q]��/�3z�f���&f�
�p���(��9��&rX��&�R�X������U�>
]�t�{�~m�rF�Ny�s��r��1+0�s�>����� �5E%���!܆��̲dRd���Y��Z����	;s���C�Y���O�P�Z��ͺ�57�<�mq ��h�E;6 *UwB�\���ՑEw=9-w�$�FQu���4�#$��pl��HK��@�,y:��e�x́q+C�%h
�8	.*���Uo���&���?\��P]܃��D)��έ��ד&c��u!����>���YZ�*����7ڢ5qV��9i\�ݳ��m��m��e��g�O���#+��/'T��F#����-���[̊Kx6E�=�q�|��]yOs�j��%=G*X���tb�DD(���j���ui�:�\������p�z���?6ѓH�5���H=�r_� f!I����H��kL����Y���6ډ�0�&�i?T��'����;�Np?=v������Tiw�]����A��l��7DN������=�.���T��/ٯIOA���1CĞ*C��.DF�?h��H�zo����&D!�]|E����çп��L�3�`�S�'�x43�[���> C;�e��0s���f!����J�~�~`I��e�L"H�YKZU~1o����j��ʌ�K�{�
0}��e� @�Ձ���MWwa^�R7��49�4h�S�-��\tQ���=��V���Ѐ]NF=ϰ��I�F<�GT�9K�G@�ɀ쬽9;W��b��T(�����1��X,쀓���V\�{��1��,�g��4�W�ƍJ�dB�}y�����'�W1��4�I�V�Q=��,�6!���b�Ak1��߈}��>�f]{}e���|n�*v0�_d��73˲K���/��������M�N�]s������{��.���S�ű��3q!���4փ��)��R�b�8�r\
��z5�D�ݑ��WW98��|_�����J�~�	�l��"�T��a�c
/����f NW[n��j�Go�%W.����p��L1��mI�_eRȪ���'M��U�$IװzQ�H�Yk�c�8�M%�u�B�,��9�KN�ϣ(�N�Ճ�'G�5#�~�߉	P�v�c����+�JG}���м�H���b_Z^vnJ���U��������~�xv�SP��ZjA%Ct�O���ɀ崹<����`4��F������R����Մ㢹�*� n.�o���i �.'�����Q~�{�?��nE�k������������}pb>�R~=u�����m�޶�P�&�p��b	a�Br*�-�/p=) �%����e����u|��ۏ�w��`��W�62�r
A[꾛̎���~�g*�TZ�9&ύQ���:�~��\=��Jg�G��G0�8�ԏ�E|$�M8���N�5D�����o�4�%�B�{.��� `}/�%*�uYT�X�\�%�]y��Ҵ���mNuu��^�hn1��+� �a\�4��"�W�d���������5���p��������I�=5'We�xY�1r�b�S��?)�����}"l8&��st�������׻��E�D�L�Է�����R�
?�2����]^��7��0�Z��ޢ��>,�~y1�D��ۤe�]r0�F0��>!%��v�Ջ����*�w��t��q/|�k�m��Ek��
>� $#�R0 |���l�!�.���
_�3e&/S�l
>"��eV��Q1m����ΪN�5b�]���D��J@rgsW7G�@�J���ydt`�/��V�_:~�+��c�q�[��lW@!8q�5�Op@p��@>P ��7aI*5K�]E�о���c���M���%�ȧ�g0R�q�\���j�o��v�*����eA��Q0Nh�Ƕ���Į�9�z��>�]a9f�S���������wn����YᣮW7w7�'5�6Ӂ�R�K���%��=�-J��i�����nL&���� ȁ���ć	���*.�[Y	aη�Hᑇ���
�	K��٪�P~���^�#8UY%��`0��:bA-2�Dd�u�#w�0�u���J�W�ه�w.
ȯ+4.��m.v��[:�}�L���<��[��]K�5���G�_��F�GN7:@�m�,�uP&{�
������m��L���g:��J��ȣ�+� �0�IҖ���}�ҋ�ݶ8ؓgVBvq�W�����wHhM�YS&~�]]}#�L�d���*���v����N��m� �dw�T�7��$k	���s��W��7Ad�(���@�K���p.x��_��qod�Z�y����mҾ�Jÿ��q'�U�f�C~��b��6V�`x5������Qw盗7 `����jQ���$��|O�gy��{��g\�;�W.*�K 'J��ύ9�HFǯq�\�v�u3���T3Z����C�ͱ�侹��s�B��"���8�L��0|��\��.�.�#���6�?���"i���mZ�d߻�_Lz1f6n�+���f@�Sە�����o�o�q�*�>�E��(�W��Yߥ6%��!��g��Bse��ٔm7���nQcP:�F.P�\v|9����m��\M��g�]G;��yE^6&-��P?hPV34R�:s �♶�-K����	��#����g�B�ǭ�ȹ�L��7틪��=�&ytgH݇�_�0����08�Ќ�*�����n,
�������Sf =�!?�����6�zvx8�}�i�K��*
�>�4hXr�]�T4{^�K�Iq����ы�k��0��ƚ�Yh�����tJ@f��e;P2��kQ��j��X���0��`��J�Ha:p�y�f�V 
&�W�����.S��{�6U�e6��o�u�l~{�x�zgRO�����?7��/!\~�Z�(��*���w|M|�)��;�ԩ/�z5Kjo6.�������ȍ�W��ݶ\�D������4���K7���:	�����"ƈ����>�|F}�A�o��T�A��y��Nv��(A���^]	�Iܐ�⤻b-W�J҇��d{������,�Ѫq���v�_�A���Q;�+]�w[����Ǚ�{�+�r�Ϟ���A_�X��V��<�����B�݀SKΥ�Ϙ4$�-�x����kh��'�Og>��`z��ϳT�j���]�dMy���|�vg�/���C�&�*tָ{����������-�g��Q	GW6G�	��0�1��ގ7�X��L����/�LS�*w�v�0->�G�l����wu�����v;����:E1����ʠ���ߜr�V<"�ǳ~%(ÑQ�6 ��X���*[�a���IC�r��� H��#K$�h��S���q�\�@
؇��W5N���L��=�qn�2?y.!���d��5�;!�����$�v�H_�g��9`�W�,�N���:�k�<V��b�v@������!�϶ ?�R�UW�G�z������4�3�'p,���"�ߦ�`�*_pj�e�9����S�xM<�	� �6��#�̜J�OZ��X��)x���T�<�UP,yl����Ǘ|�+�Q�-�C�.�9�|�� ؃���x�#�:m��fWJ2���� &6��:�lD��E�D$(���C���q���$2����(C�[��7�F@����/�*�X<�q�3<�e�/���R`�;]t��u{ѯ��ăwP�SRq�@��@������.���R0ہ�:!7�G0��ڔ�ilˊC9� �/}XPj�"7MS5u"�Rn�f����r,6�����d)6��#?Mp�E��~�bL�P��<�����=�����v�/˿ͯ�wy��`�[�A���%C���OW��_��k�s�x^��|��f�O�m��G\��HҙxkU��еi��O��f����b$�,K����,q��j4N���b4U��+m�_��s��"p̉PU�^�D�\�8b��ǭ��wܛd�(jzu��`n�Ի�_g;˩���Ns�ӓ�o���y�{�]嘬���|�%m"��v��]�.E6Ff�h�w�83Hf\Q�f��H�U��j�PT*�@˟���$�r"\�g8lOუ �'�`��A)��hر�⺕?<��*:�����������Ѱ<��z�~�ŏ�Ctx�4��oK� ��1�c�u�t`/�ٞ%K�"d�GT�L	/��KT}�8�7�*�
�M����V�1g.�P�,g������+��c/���z�����]$�[�_���u��O�>��EG	��A��M�� @����(�I����m��6�'��0�>J�3���1�m����j`�j��Fne����!� )4 - �=zլnX�h�|�z��@c_ɑ�d'��Z��_2����:��w�[��kź7��LWɇy�X}���Wb�E����T���V�fz�z[#��F׀c)��������[w1.T��n$�?��k�����Q�C���<Lh�c�L��#�@�~/>��m'���2=�Z#��P��k�o@E��/�ly|J��@�bUILU��E&f�vk�<�å��"`Q�葎��GQUHMOg���NN�F�b#((�t(m 	MqS娾����8ƾ��)}������]M#�	9�R��6��[u�Ϛ�ga9�%-ڨN��pD9!�IuIr�˕#;�ů	&b�AĀ��/y��c\�Հ��~�@N����gXlxVHYEB    c945    1240\�6��yerW�f0����Μ� E �8������j<�U=UX��b07PW.��
��|1�ƘI{[��<�Ҹ�YɺPO.Ih�C�. 4���;Jc'�ǲ�%ַ�FT�K`�y���-�h�8�z�Jؽ�7)�Xn��A9��p(�Zv��$0��岇+�k�OZ8�(GY}G�0���8]^����ȵ��m#�zBaHB䰣|�N���9�Zx������-닞���i|�k�!P��ڱ��
/�,T��dA���FЙyÍ�&�f������o�tiF��{�{v��xY깑Ea?����t��7�i���\�]�4Q�3��M��TgDw$Z	�/��WQ˧�ei��*o�5i=��Ebˡ���a�,f��c�ӯ�ٯ�T�^	}�S0X�2�-�W�=%^��5�����7�ew������l�P��F �V����,
��eA��L)���X��A�zD8J���L)�QoDl�K���J�d^G\���:ݺ�!��`���8���Z1Y�>$��x$���Kނ���"���>���8+�ê]�L�H����=�/��K�c[6�X߬�p�.�xP�kn�sU�p b��aą�X��V�����]��|U��ȸ���9�߇L�qA:c��%�P��\�ɪ3%rh|�IGP�p<[�a�
�*�E�!K��hWl�
t�7=��d����� �2���~GLr��z��;Q�[g��6����5.�k��H�k�/�N��)�z��
��B�j�O<�ES�= �q6���=7s���e��u� �ube�Q����܉G�K������.t��N�IR �c��N�̀Ę�������dG,��.�!�§���� z
Ӊ�9q��$�bYX�h�����m�O������b��k�ux�Wv�x�?y���N��%��V@"\uȸ�N���9�<��:�Q�0f�mO��8���F��Y�i����kG���Ѥ�L����uI���PK
�&�l���Ԑa��xZ�R�-�Y-wcd <p�N>��t��k��$pk�������O��)�@o�n�tn��*����ɪ"�h�o�Td�3W��\�	#P���">���;�;�s���੯��&�ey�^]/A�k���O��'��2��]�zl�j��]��&���A�[�뛔Bi^�7�Y�9�d�@�'1p��A��:���he��ڄ�QU��~����)�"-����C~~��'=�����|�p��K�3Qڲh���o��p���%i:����:�`��aZ��OS�j/����t뒄��xB�����턁?rj��NeF#)~�� �I�"�6�q;��s&��Ҷ�sk��_.0�# ��ho�]�F$�,�v������'�I%l+�l(���l�y��G��	�D��������
�̓��V��I�Bj�ؘ.$ǥ?�H�7ޕi�c�P�_�9Hp -{.	;���;�}@a�s�/Q����f��4��1�e+f����*�ZD/�|f\\*Gw7���j�7��)�g��k~kr����C�5�T����ʏ�W$6�&<�W�5ve�zkTI1�����WܒK�u�W@N¦*�'Ini�K⠉�#�4Ȩ��8��}\�+�곩ewf���z�����g�~�����$uKB|�
թOC�?�Z��k1����b����P_�W��ҕВE����B�J�?2H:���K����,C�4
�+��=�=-c;[�`�����˞ֳ1�.����!%������b*s�b�
���z�v�����j�7m��2�^p�ElYR�Akx��kQ���^Uf�Y��?�8
効���Ϋ!��T`ߙߵ话0��]%��{�ʍ!Z�٣� ��o�x���x��2�Od�d�Cvy���{�$4�xRu�U0����x��V�L\pc��M��Dj�L�޽{y$�0QSVᇫ9�K����I�-�.$YȲ��#����)���Z�w}n����)=����e��db6(xU�-��EE�ؗ�n���7��l��f�U���$����a��K0�*1�A�/��G��Ǩon`�8ݳ�&��Q�$�욁�4���!�p���Mj�zo������>kƞ(`E�!&t�'(�NC%!\�ڬ��j^�n�b��gU'��h�Ɔ��$���2:"�y��X���WgP
G&�D�*>A@�����[9Z��R�:P����J%��I&�e5�qH����O��.H����xo��C���r��T���I�re���e�f>����b�l;���7�\�W�֖`����>��8���R��-�Y�?�$�j�Ȑ�*p�Uv�*��F����B1k�����lv�JMSk����7�����|�i�T���"1hj"D�o���TJ���iflP+~ƀK�h4��g��6��J>�d�I1@�dhkƎ��	�}W�"���R���A�7A�,�١�_��4���*݈A�k㭎
���������{�-�5���1��Ή|������Tж�^"������K�L�������,Jy��L`�Vmv�e�&�^�f��0%w[h�+����)���>.�~�����M�cX<�Z�InY�H'Dy��6\D�;qw�� !;])t��S/l�:�J�D94�}�Gݿ��&���M�~��$�ԩ�o����*��{��o�����Z��p��4Py^c�����>� hZ�����T�b�
1z�J�|1iF�X �:�R?�IW\�Ĺ�B�c�~����H]L���,��2��c�W'�`	����Yyg�hF�e"`���#!Xr��ů�sݛ�n-��T�i_d���W�8�����z%��s�3��%`��C
Y�@��Up0�wG.^�^ 1l�I���ҡĠ��j��s���d�7^ʮ���g.����Wv�|Ҙ�,�9}�og�bv��P5Oh[n}dL�rm�*�sb\q�����2�ƚ���b�6zE��i�q�7ȁ�����P΁�[��@�T�&��NUT���}���?�������
U�ri�B��u;�f�FR&����ax���ya�%�S��i�jAO�eD
Bu��uzo��v��1���`��Q[jH�!�D���a�#ڨ�T;�aJ�A��Q@����?�p�+/�eM_�Do��߈[�}x�ү��9Qm*=��Y��d�_G�Y�*��'��͚�(�F��s��{X</�猪�����Ɏ��gl�LF�֎�ɞ2L���(�+����jt�&~�Nj���T��S���9�Y$}��l��C�!�c� �$2�e約`�r�'��J�G2܋d����s��.���Q��Ef���'��E�fN���1>��^���z5{�P��L�;�?��{#d�1��u�#�Ok_�޿�[eXw���A��jdF�eQBgj���ӵm�pYJz��	sB,m�kg����n3Φ�z��x| -�h=Nϵz��gm=v#j�q�W��b��O��D�լ�IH����:�5��ذee���Q���	8݊h~�F��
��&W�!�S3+Q�J�UܵRC�~0�F�AɈ}��\N�舵�K�T��j�=ad@
o�4�N��ӗa�{�:d�4�-��<N�P؊)={*DʺQ�_��>
��#k���
�.�3�MS_Z�i��ai�7湉�f�K�A����*m�����ePJ�0ʬ��'��$�\W�*���A$�Xu�oo��y<�L�v�~:-�oF'x�M_���f��j��]�0�g�rE����Sl�^����1�53B�:M�!����W�95����=��}�9���J$Q3'uK��Ȭ��z�R�)���2y�|���=W�d�/�FGJ���ć��-U�Wa���$��nN��u�S�=�/�^�LM���8�Ⱦ;v4��&�k뺣��?S�yq}����$0(�\M�7KH��L�Hm;N��<Z]߄spa�J�Ӈ���Sq�le��9ƺ��l-"m����35NF�w9����۠���dH��i
�2��K����.W!5��:VG��Id�Tף��&�oF���` ?v6�_0�\����KR	����y�'��%��wl�"�$wE�'$\L[��͂[iy.b*�b&��|-�&QF�#�1Jo,S��}q�7�+q�^��H�V����p�k�6m���B����C*Чo�`�'�?E\����Rh�����9T�eA��J������&��WӢ�}�u��j��>> 0+ҴS䚬�g);CL/| ���
��z�+g-!=�~8�BrCY�EO������ĭ��N[q�N�K��e�sa�>_\�?�!Dq��O��G�$fj�Hp�!�`���5������8+I��Z�7�}� VW8>�I����grlo�l�F����z�u�^�i�'���-2��2bg��{r��_��~�|n�N�.i�|cYQ�E_y�/�+��|���u��3�vV�9>
xr�v3�.�*��X`�Z��#�B�,����Y���Э���Ϛ����,hx���	L$f	(���"�HE�5��Z�7�"7�[��S��(Ǣ�Z��og� �����}涅��t