XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:Y��D8������}"�7M����I��!�[bǹҵ}���ț0I����4T�Rc��p��4=9�H����ak.s�K��TeH��<�nXB��ڥ��Q���S[���}�������%@�6A-h��q�,e��QZx˺�f��ݯp���M�1��?�b��!��-&# 93����VZ)��w~O�$1�����VoiL�9۟�On)G	/����yY������f��:g���(�p{8��T(��!)�-��3f*[p#�I�d{���AE�9t􆗿֗��#+(v�q=~ɞ1�_BJZ�T�R�{ͅ�tt`��@��`h؜�L�Q��L�?m�$�W@k%�!;E�ɪ�6��+!��Q-Lw��-����W�lT��#�,;n.U2!�)/��0_��a�FFO	�i�3�i�����=��͡Iu
�;�
�X�_m�R��:�V�_�����t��3���h!�0������xc����E���������27,&��	T�fr�_B� b�Z�5J(ѴY�?Ý�ٍݖ��_�I���{���Z��zه����A�Kl�bV���ìj�E�q�������/^�.A�����b�ϥm���	�-�p��p^b���I�_������g{�f�F�wx�2Sc4�D-��7�0�
@�/F��	�D�'�Rr��Cr��"�$���P�D�~p�8@S�B���5� S:�~{^�����|H��pf�败��oXlxVHYEB    5d54    14e0���zߨ0�3��CM��?�!�O
��H�ᡭ����}C�M���D|6�/ >Z���=ʸN�޹���:����{�jh�S�j6��=�{����4G��v�Z\���D�{�ㅜ���9B�~L�/�O�8ɝV�ȋ�rՑ���1!7�ʬ���4v�`�s��S�"��MKFSϞIr�S�\s���C�wl:�v�pWJ�1O>�̡��ω��J��q��n9���OD�$��ڇ�����|~elI蜣Wؼ3�Z2u�̠�f|�x1˩Lk�Xhi�ovr�U"����E���	�bh�-���o،c�����LT���E1�O
�u4y�;�<�{�~iZ�c'z]��C���U�*z(��W�8��>�)��:kM�0�(�w��GF
>�����ϏP+�ނd����b��;�6I��;?���F6���5(�xpm�ۤ���*e�
b� ��Թ����ݰV��������Ǜ��z�F�3��!�ԯ�IT� ��zeɼ�z�sn�N�z����H�5�G�o�9��� գ��ÿ �q�sa�#x� ��)�s��݀��?1%R +Q�\da/�R &���_~���JQiYX�4�%��4R-�'e�idlpa��Ȩ7r���`EJ'r���zh���q|�� /�n�[�-��6|;r�t��o��l��F�n��S��,�g�J�d(���}�D��?ѫK.�O� A��ã|8��k��4]���Z����(\)�7�ʜ͐/�k�^���B�pv�h�8ߗ�¸Jh�������I �TZ��n�/�Z#���7/Na*����%j���ҹ�b�Zd��"E�{���\y�-X���O��/H��Ϙ.<�ˑ����N�}X������$�|z�pmo�� ���Z���mk�#��v%^����.qJ)e�L�Y��l����Q��͒����_7������F�˒�7�����<��٘�Z_�&Hm_�^�Ǧ"��G*�hk���t���72�!�e�_O� #����Mᨋ��R�,�^���i�}uU	���NOm���_��wgR#�&��P�y���z\����K+��'
��������(܆%��	�Z�m��o_b��8�ӳ�j��V�oe�$��q_�D�u�^���]�4�e(;�e�e׈�?9E���ZU֨u��j%�wVC��#5�i�?�����!�{.�����L1��"Q�@`Y	�]K�m=�Z��|;�M2��G���H�gh,��n6@�`|��,'tBy�Q�̌���!R�O�%>���R(2���B������z i��:�7<q�c`_��{sk�f@9/ ���<{mP�ŭ�I$H@��e	P����Kw��o��z W�	�\�|@���l5 eJ{;A=���d�#��u���t�K3ULO�ƶq
4<އ���ΟB+�������R,���_J�������������	.{ꍇ��o�R�k���q�6/�z~�?�w�5`�2�#ZTY	0*�L���%|8��Z����;uK���j�lqoJ�<��rH��ۓq[�dbs{�b}�-����k1��/U��]ya 9�Av��� �l����������Q���%�2"�Y��rhR�@ \�ᔵ�k��Gx��تʆ�a��w+C[����.���'t�|:������a����_6�",�#�g7���|��s#��K��4��$eR���?lb�7�������{��\�Sz�O(��jX�����Ţg���{҂8h]������u*eZ��!�3��$#�=F�!C~�l�0�b�J�]���T-�tqtW_B�g�wZ�A�wZ��D�N�<.��l�a+�	��g�w[ݩ���l�;���:PN��) {�=��ȱ�o+�A�n��QXaor�o:S}"s�6�Fv�G���Э�\���#S��oU�`�*�6�µ�  ��	4E{��BOM�-����
����B}�>���bѣR:�s배aFޝԩ��j0I���y�_?1GJ�����B�,����u�e}z���������Z� �X2dkT��k-�"�*V\�#��س��:}��|{��_6�a�VDhO�:���C��pd~Z8�41?r��M�0~L��UK(���p3�*s�mTZ<�U���&����#n$M)��[iO��-*y�ʳ�Ș<p��w�(> ������l�B봂�����yjC4�Llnk7��1���5���ߺ��E�C�	�>����Hh�0S���K������B��������Lap�=��C�.�fP��on��z0Os˙8zj��2ެ����Gz{hW oo95��Eѧ'y>;�<+��5lr����3f"5�Mj�^[���0*�w��
�g��7��э����`�R}Is\�f����T�ҹ�ܗc��	�vNNU��O��R9���?�\t�A�3��#u�O��Wj��S�6ܸ�q���9�(%	Rx|uߞ�W�5��!.�y]���u	���^e��W�Yl�L��ӜA�?�<�r՜��;� T�N=EYѱ{~ֶ�=����cI{�}��z���69��u�e�k��X���A�J9��1�C8&���Y����w�a�T�;�{u��Y��v�^~�����N�p8!|�m6y�]u'N$�8��N�ǤX�^<��92�h�"O�fQ���{ݎ���!�"u5�o����6���Xc4��d�e��Jz���t�,�P�Q˾{�yߗ�,��q��)n���ugY��lغ�r9NĭGV��6�����bF�K�����JёΦf�;�T#�'�x��.w����P�-Z�����5�H�n3!��k2��j�V~/��K�m[�Yb=�_��O��h�L�xCf]�Ź�� '%hA[Sy?�X���<�(�y*�%������H����Ԥ)I���ҍj.�A#��Y^�����p=���HG��b��K�ڰ���/=_�.6t��)�ͷ[��8x;��׆�Am��G�W��Mhr2˞l%�9m��&���I��Ϋ����-�ф�.}�~k+�l��n�`�yF�zЧ;a�)����z�Z�ڇs�6������Ӹ�0� ���zV�n�4d�
.�~�
�g�"|]̓y�#64�[LSщgy�g��~��>��R!�n?�
�'���s����|_D��4L�L�w�˵�_i��R��-���z\��~��U��N���f#z�
V4�B�c/)5������s¨��{橙q�M�0��*t,�Y������=��c�a�u%�?�~�!�/[�
	P�K�]s:Z����*:k�u;�VG;�v�U��+~�� ?�)��7r2��P�A��嗍jkNU}1Sbk�}�ne�^���a>k5�*,���7�ͼ�?����}��tO������Er7:��z<�pI���g�lջ|ۢؾo�$�y��+�U�+��ߥ�, ��" y-�A�WC�9O�ҁ���%.��b	ܘ���Ra�`w<����_�5������]���P롤#1�	��5gZ僻��X��C~�C��m9bA{y��
�]y������j9�A4gP3�ӟmtC�Ut�x��%n�4h�t5���I���]����ϒJ��asA*��`\$��~j����D�E��2V�8\�֥�5�I��ch����Kei� Xw(��\�I���G���*�'���H]�OFy�u�!�m��/o�%� ���~����\Ǽr��	;}-��~H���~�!�n�|~�E>��35_��e����xb�
�&U'���}�:���s�/	x5jf����9��jQ�ނ�q�1P3�R7�As��|(�z�&�KR��/��%��'O怊�H6N�T��J+�tl	���,���z�R���U#�D��ۍ���| ���9�J��r�i�/!��٪���ek���V��t��W��dhl1^\���.�����AFR��3��;�N�+���כ1��f��#*��aM��	X�ga��'�R\����I,���|,�3۪jGSa$��_+pM�Z*߄�"��@�?L��T4��h��WGF�Z0r���!���I�x�%��z�7� #����:e|���0�mL���~�OF_�В�s�C,n<��r��P�g�17�ബ5�eD�cX�tS��s�w�]G��^��}�I���M=Z	��	�Z':Y˝(�E��V�.���><�(��p����0&82A�ʻQ��ilh�YH����*�gV�,=��V����E40�@ca0�$��iڇ���w��}�$7:N�8����;���ʿ�ʄK�n{�&7e `�v��`F�l,���t����È+� LϮ����0��2��v�c�Dh~\S�A�r˼k߭�}�Ř���O��ߵ�l+#���^��dhT�[�}�U��D,�a)F����pl�m'�B@#���N������ys��?\�cjQ�oZ����X
�+O� vR!e��d;���=C���%�*���?T1̡Qx���	jl#�� j��閗�[ߩJ�?d:��,����R��������t�F��S�h��7(L>��o|�є|~7#�ڟ�󊓊Q5��}�4��sP���]��o�����i!�:"ej�SC$<iU���;�jkvl�*a�h�c��NsN����a;�]j
�og�ap�w�pZ���\?�%�l����6�W�Z���������C�#��zQ�S|D-������*�� XP�+\�����ґ����ߩ_���ҝ'��6a�'|'I#G��y5Ϙ0;f�}"m&+i�`2&6f�@V��U���qJ^��Dr��S����@4�)�l�<��)1Vf�&��J�������yy@��V���}��:�ج��,:f�R����� MӍN�dv]<q�J$�W�������A�ĕ<I��˂���p�?�v���Z���UA����Z�2Hŋ����jV[6��j �R)���y(��ˤA�'>k��b����_B�19��gJ�G"�H�_�s�x��1�5���4_�#h����״� w��>A��~�b��ʉ�Q�0�B���0K1+��O�m9�k�h�J!E�bN���P��1s'�b�j���b�4�o�5�R���\��Q$��+m|B>�0�reؽ�;�'wIV���V����R�!�]�݉�����8���ɒu��"N���1��=��