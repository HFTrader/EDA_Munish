XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������^�56
����E��U-�#k��� �L}��;��hӿ�l$+Ȭmj�_�,:g�E_fA4B���ڰ�2O�}����
q��2�3��y���ݤ��p£�T4�J��30�Ά����ɮK�@\O�v���~@��	�)^���,��9���$�I �Rz�l�b'?�$� �Ç��JA[�������&�m�NW��t��~u����!;;1(R4�3�M^Y�.�0�7��{?P����ᦸRMG�ȼ!�6a�''�[�ɢ�R���*��#6�4}���Ր S�.4gTݱR%�I�(��*h�����aIl�o��bo�e�D�2��� ���~09�)s0b��N�ӹ�'�S2�9���Ar�B���BN�o���6Mڞ<FF��%n��A.����>q$K��p��}e�q����2�W����
�ĺ<�0B۔�&�S�.�������d���o��B�����[������%g���+���.�/�|^kD��
�`�n/6�0ڌ>�4U��E�	��X1����d!~Ǻ�W,N?ciT�V�ԧ�� ��O[U�
���C��O���5���xB��-8>wK'�ڭ�7��\zQk��抶 ���z_;�22�
BmH[$�'�O��E��`*�V:9{q�)�#�T7Z.�W��'���F�s.�#�Q���0��Y��ch�m
�<�&=��Ȗ���j�WPǜ�1���'���-��WB�����sP�
����G	�nXlxVHYEB    8990    1bc0��o��c
w5P^�w�4h�ّp��VSS��9���]Rʧ�Mz��3�Yv����eԋ#�\8r�����k� ��Ƒ�҃V�;�7�O�a^���>�a'�E�-�+����98�&(���ջbK1�}�W�C<����$�=�W�4<Z�;b�Pz{T���A�G����+�y��y=�
�h�k}#g�d�.)�/��A�N����D[���/���X�i+��t�׫�@�4�ľR�OhkPV-e��}E��w7�]��<���R�4���T�j�YZ�<G��|�(϶�9ވ�--��7����ƌ��QH/�ם]�%&�iF���:i�U�')���5�y�:��~5�]�M���A��mGX]�p��䜿j� ��k�����g�(���̫�n%F���7�3=��=���t���h`Vb��ZH@C�dPGGy:��FbK���.$��ՠL��FDl+�n���$�4��L�/X�h��و'q
� ���Va#���q6v�&���$�ί�I���f�t!���4j��g_�x!��!�%)'L��M�0�V���M![��� Kߟ�ƛMz���|�Vsf�&�%N`�yq�G�,`��.hFj}!yc"��2�<��s�fEZ�]l�ez��O�-�`Uӽ�n��!�jm)�}v���|1�̭����s	F�m�^�!"ims��-+3@hL��ΌU0�����\N��P9wE�h�oI�%��䮧�Q��7O����k]��zhU����E�gzj�����i@����1p�|��W�.j�<���ޟ�ؖ[�'[Pc�l���n�[j!�QB��)ehȴ%k��^p��"d��y��FCY'�6��F�|�x�k�r_�����DL/�T`�=4���u�M�� ��t.�_H��al�~��4��樆N�N�kB6S,����w�/q��c[��z�g�V����S�>4�a���B�{�K�~��(���D��z@��]-�{���
����R�0�ijI=�8��lMo���`V����*��٤-�V 2��5�Z7�N��	ͬ�y����G�o�2/-F��W%0��O)4�Z�������J+��z��48�Ӷ����:����<R�2i�V�?�,yF6[X�t|�U]��^"�u�Wb���j��E���/*x��´\�E��pNر9%M��i�l@;������y�tdI{���f=ۻ�`,q?�Q�j��FS��l���2�
���x��sZ�}*L���7*����J>��wZӜ�Q&�({���	;ȷW��" (�a��jU�E�R��I��$�Ju�Ǚq����j�}\:�k �JI�����3�{;�u�B�D�-KJ�
��Ȇ ?����Δeڂr�)���T�l_|�#����(I�����p�	7�",WB*}����}����^���#�F��(	7 �ysɍ{A� �o��U� |td��hw@v[pZ�3��Q���Q�k~�9 ��L�'��{j�T���buQ��s������դ6�A%
Q��2���GǺu�Ǒ9qx���= �V)Eb� \����%���L�8��,� ����{X��cL0�{�>� ��,3]������_�^6m�×�� �dX���P{�R ���1%�������v�F����C�˱���c5��n��\"}���'Ñ�{�s=��ւ���!o1G����G]u�y�����iEڴ+,&K��T��	��t<���SDX��A��m��0�%V7\���%a�9"�Y���8�$�/>n����_f��?K����n�C�T���һ�q�}y��¢#��8�P�l�-������t�4QȽ!��&��;[	n��v���i_�g�ͽ���&�!�2��c�2Sh����F8�9T�p��1+��G��1(�!%\���dp�\9�&��ƬmB:�H��ؖ�������n�1b�1]Ԝ�� ��(�śW�	\7�q}]3o��R����HS��'��*�����9�X�o0�1+O���[�В�}K'Z���kӶ�da�b�v�[_�,`�������8;�����G���ܼ�7Nć��xM���%�;��sa8�j��S��M��3�� ����
8����a���q���p������V�孵6��R�����l�9���ά�o���GI�J�o�"�T5��Y*��<�4��ҙ��A��֔��!a}���{�c8��~ž�mY���G��	�g�y�Ͳ�ʠfl�v�dk���΅Ҋ�ǴZ����8����PT�M��|:�o�&w U����2�M�d�@��'&{B��-R,��,�t���0<n-��;jB���.(`�������I�M�Xd ����3!ܬ�~�a˦F����o,��idWtl3s＞r�<G�l�|���R�[���;Q� ���� ��a �1:U��}Nu�{'�\�n����-�]�r�=/�V)��~�]Nۍ~?��- �����%��g$.�?u9�\4?�_m�̴�ގ�gC�4��9��!�I��\�{jޘ�Z�����-�-behj@f�����\�G��*�]�U�	���lsퟷ��ư&B�=9��lЦ����� "�k?��!��Z�r/��Ŷ��g�$zȦ�J`������:�J�	T_"����`gC�Xx�~c�)N��Ez����]��9�sLQ�����e,��x$�v�D��L��ُȃ+�`[Ʌa5�j��{!=6u��	�!��OS��,��l��a�
,��z�?��Zo�*^I�|ZJ���u���g�6��en����6�3���3E���*�X�C2	~}��䎨Ts��(�*2��&�����JuO?A��gh�5�{��]Y�=�0�Х�gEw�Ȉ�E���؟�����;׸�Q�V�)UN�?�&R��96S�l	�4L0�gf�z&r6J{ks;��-JZ�|��Z�P}���bj*��?N���R6�c"�"�dP�Q��&J�/�#%#���T��C7�i�m�7�p�KȲ=����1�z�Kɡ���=�#|��p���0��X�B��i��hv;��&���[�*���� t��	�/��<�'+Y`N��m�M�Fg�*�K�SW�Mo�Q�]�J��8�1th՚۵!�!u�D��ܱ����659zDo�w������K@�[�Y�J����8=a[Z2�j���L�G@40�hB� M@�w8f��*P�$�*o�z��;As���б��CW��U��&P0_�
���ms�5��Wɤ�"�v3��2������ZM�V.LT���y�$�Sȷ@�4)T19)�Tx���>v�=��u�s.��VT�v�����]#��c㪄��GW%e��+���x 3��}"@��nS��7����h'Z�Զ٦�k��Y�U������b�2sl��v2�zG���כ�Z(2\Y�AK bB�H���A�b��n���D�� Q�������i��vޒ�c=aϗ!��%(ND����zsɀ�,�I���a2�J����j>�1�R��?m�|�L�ӊo����XY<OI�R�j�ZN�"A��Ԡg��ܻ�$��Q9��Yΰ�?�6���Y+Q�70E[����G�� �m`]��XuB:[�]u�%��v�%Ԃ�l��*ƞ��";(��"��0i�n?�Kt��(w�@B���H��M3�cc+=�w�C!n��B�� ���$�(Ge��Q�����K�������[v{L&Z-���G�$����4����m�ӈ3.���7�9�\�~.�V�D�L����1|��ʺ*���n�21@5��}.�{�p+��d�<)�͍M|>�"5��^��_mP�%�+����A��I�u�*Zj��Ѥ��\�"S���BO![H\+	A^�&��:�[�O÷z������$�АZ���O{��i����'�(�%�~�ߖ-�ٻf���B�6HӊV���.�;zI�7���$JL�l$(G_`�I'r��$2!T4lj*w�(۳E'��5`��{�7�3�(�jچ��WG����T6�8�g	2��Z�*�g�3Abd���\��o�������S[1/� {����%�Yxc�1�3�Y�y<E"\@���̵�;W��].�}��]��\e÷(>kK�J�K�#�޴,[����_�9gA�5u�@��r��X�=�I��q��J�0@M)����)�|�>��%×�rdo\gQ;���1o4�o!1��Kc����=��Ǖ�,��i)w�)L��D�0t��˫��*�Z�

5������'�4��1-�&a3��.��5���+0�	�pT��Ļi%�������=��\V�z\,e���� ݙ�a���(����{�
n�?M��,?6 ��g�m��|�����������A�#}���"�VA�[�y��v
��������]S��4R�b5O"J�Gi������NqU�F>鿄]R��F��k�����X�H���A�ҫ����=�Eq�8w]-������S\*��.e� �P�p>+o����������uZ�w$a<F0A1<�	'��C~���p��ل�r�Z0��JD0E]��[��5��{�����^?�1�r����'�WEG96�} y��U�=B�����P�sͥqS֭�Զ��� ��˼���~�i���ޮ��.��v%w��tv��4W��1�Ζ��1�ۉJv��WV�S�="m���	O�TOZ8�K�z�0 ]
���� �+�����$W�����2T(����x�)�~g(.�2ua=;Φ�#�Ωq��ML ��9��^�B�!�s�J��Ss"�u�-�B�c���	mc�PX�7�c����@�N�m�)���>�a�~���S-���!�,��eyT��#��o^��DTW?F♰����LY�����  |�S���p�w�D�Ο��K�)tO�_2����+��iJ�줅Ӏ<��I�9oW�9���6_^�Ɣz͞��9�i� /�{Q��w���y�M������X=~�2#���'ޯ��(�h���nv]�:-���N]^)9�^$-Q�d�B�@ڮ��\����n{��V����)X�ѪB�܇�=6 j�,��)�hge@ �@�ӊ'���P:�"������M����ŭ�
�؈=�>�.4��DW��;(R��S2�;d>�CP�T���whb7Ϧ�`}�F�S@f�x�6���e�`���%a25��b����V���,6��S~}�Z})uu�⑖�BP^��:�/V����鵂<d���=gp��S���$��Ax�b�B �Ӂ_�2�zE�4�2�I�#q��vB􍬧�X��ȽMR������E�Hnº/��[8FҠ�o7�Lz�јlWF�AS�1�٦����a���)Ŷ�~�<�j�R�D���`��A��}�N��Oú{��0���'˖_��H�1�mk��� 	3�k8�|QL�^d��W{��xҳaAcP%$e.�C]<S�L��Ks�<Y B��R1�ӟ����x�ga�9��;I��[�A����K>Őkr� �W��l�せ�;F��\y��e��~ɪ�Y3Bkb?p'w�ZG#�f-�j������Cx��}o�T��V�+ "�+M�'��|� ��7;�"���x�PJ(�t7�B?�~zY�=��
��#���)JR˻��ci�)��xpJ]��QD�Ϩt�����b�4���me��;���x�Ǜõ�h��݂�%�ʞ�[��L���mpA���SX�]?�7
�D�;��D���0DQ��yI�}u �;+�oDM��J�<U�r���/�g�Vf��.�m�@h�T� �����lPC�,{��������0T�
d�����p�N�7w��/��1w�#�Ldz�j���9)����a����aD?'@Z����g#y��-99[+��5�r�_X]uI�5���
I#��y�����q/�����*����l)�$R2L�!t��R;�T
���w
�Y��d�b3�"u���0]�&�揇�7�ëe{�N#k}�a�����k��ٍY$W��O���C��r9C������>Zه4�� zR�"���2�g�5���/���O���θ��H�'���AYieT(A�D�`q��uV�� #L��;�{\7���6á��r��̄5?D�)z�#-,չha>0��>��s?z�I�*@��N}G�;�L�-_��՟6,���w}#��o�o-���~8�(~�uZK�P#�@L�N(yR9C���8p��qJ���c�H;?���c��U_"G�@� 6E_�Lx�P-�ٸk��pʭ��m7��Z�+�3"��ɢk62�RY�R��R�ǻ�������t��\?gv�-�5(YWʬ�"��n0���.��+��:�u�e�UK��5���9p��Y��1�ndV�iB�դ�����{?�ZQ����T�K��*��p���M;GjFwg���+4�������3�*�1��)�Hs�zBi�:�59�x1��/��:�D��a8�>T��c��[D����#��D{L-�^m�9����W���P74�RYB�9�9���V��ɸ��g���e��&��8]~J���^G�a�C�3�]zTX�x�?Us�y>:.M�� bN��Fx+ݜ2Ē��:p�S�':��k��H�������́�Z"\V�O5�R����v��������k)j���'�s_�G�R��Y1C ������&��F�L==�t��D��kc�9�1���t��y�"Q�!�$t%�V����U%q��㝓}*%���e��V-��J�@���K����E�r��[���xɢ����S�b��h�|=��c�~N��ܶ��VorAl�?��2��:��G�7��*����"��p���n"�^�p�f:�ڕu�ŷ6ѹ�]Q�nSh7c�[Zk/�Xz2LJi�i�w\����z$����/�`�}���+��o#Bj�ř�z