XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����yT�iN����mS�s�@J~�r�k�E�LQ%F���~��h$��s)�T 9��7U�%o}�����<�[��U�k�o���Ŧ�BB���\#4��?���U�q»a������q���?�����Ӯ6K�M]H�oia��GW`D��{�l7 Kg��r�"S�m}���N@���w@�0勪�k�j��9�����a���D��@�ڱ3�w�]،^8w}D͹�Z�9>���w�9�hH
�7g ȁ�o'@�%��V�/�e6DRK	���|Kc����$[�"�^h/c+w��U[�"�g��Q�X���J��t�^�4�+��B8�:�������m\�^��FtJZc ���V0��4U	ƦLS�_��\`���3<9��U��u�����bj�a�c�����@�Kj����oy*^�5���[CRsZ�&�]Ow�*����}��@ق0P@��6�-�,O���Le��c�q��٬���kr���l�W���aa3���K&;�W���(2Ɣ����~E��9�.�?'��Y �>h4%B�K���9w�c�Q|�jҐ��V��x}��N��K�h��ˑ���~)/�����kI�dR`��>r��?'��Ō�h��t��̀]�,�}k�΅LT�`�	[����LM�J���@R��܃����\��&^~���I[�r���P@i3�2	 'G���Yܑ�1([Ͼ"�n|�5�{?p���V9�R�����LЀ�^��=��XlxVHYEB    7744    1780��8����w2P�jk �̙NROkH�ifI���,Wq ��|aA͢���5�^���l�@5R�uE�#�u�	'�[�3�^�
.�����.��֡+���+0ճ��N�D����r���]��y�ý�C���8�}f�qj#�^dw�S�1�q~��_j��
���#��P����$����m9P�RM�8|&c����mi�6G�.�������ǖ���	Q�+��.�*���x��7�X��Np��+��޿w��3��p����~(5Z�ȗp8�S��������
f/�V� �������aT<+�HJx���)'�΋�L�u��L=
����ϻϜ('�bc� ^��)�5���{��*���;��6x7��@���￙Q-�p�� �� g��|m��]Ni�3:�oTf�8dmDU�W5�-��x�&�m3/���������#&^���.���O"�E�%o\����@� ��G�a��'3���Kơ�:�*�j��~����˭\W�V���K�u���d ���i"5���o]�eΩ?�=	k-����/"�]�vA�" ���[i!ȭ��j$���oه�U�<��ߨg0m�d����c�ߔ����o&D�C9R��؝��	���ŵ�
۳�������*/�h(�#h�a��4S�%rH\��r�=��]:��Z[;,`jW�\8o/Pp+�5k1>xT���4��+H����W3��[�F��$KLw��F����&DC�\���7ίs�@k�#�N�w�bV�T(��>�v���?���F������!o(_}3��m��11TH��Z�����Gc��qY/�	�wC�^)�e�)��RI�e��Y�M�].��3�8�Üi<�DN�S���^.Ţ��'�HA�(t�y�n��]	�j*�?&���m�`\e�^��3L��+��d�n�e���Xo	���-"�W�0�}�@n +m~y�{�	���ע�/�y��H��V�ڽ<�d��{�7](����Ç������B�*���&}c��}:ʝV��%Qɜ�{�chlO�x�XRc3ȔmiƉO6$	?�U^��
�Ն�ْ��"ڄ[�7qM3��VJ1(��>��X*�
�N��qG�6ܨW`\z�b��V���Kg�#��
xKT�c����V���S�	L��ɳ̻M��{���|`WG8���`������#��	^?K��H���~���E�Et�� oo�\�E��7f*۪�
�F�`( ً/��1��� 'Z�	�ܾ�٣\n�q��y{<��M�N�?�yY��A��閳S[ym��"�D��%�"wݨ÷A�k� ��9D���n<��_�;�Jq�?Ot=:a�PY�Me��DaCU�!Ϝ���v���̵��E�LRI��j�w�b�7��"2Lw>nZƩƊ��NLԯ&5�3��`B/��	�$��t�RVx��K�`Scke9�ˤ ��:�N���.�xG�'�X5R���OTx�m>�UhH�b�����P�	
pۤx�;�G&��7�O��f)k^`z3@V��sc�>X��\]���%b[�OP�,�lC�Hvk��2�ܧ��$"3M��<�����U�!j�Tn6	ᴯ���ϲ�Jݠ]"���"�ʔ��9���&�"��Q>	�[���c�
{2�2Bޒ{d9.Rt�� "m�vG&�2�)}K@��%����ބQ.���۠>DT�g���[?���0�����s��l�2ߨ�]P��D)4�y噬`�� ��c*?� ����9��]v^�X���b(��kƅ��3�+����U�*�!���FmT�0O�n1ꇬy�f�r���DwJy�lnM$�+�83�)_z��n�Џ@؄�E;��>��"�	�97С��*�k��z�^*@���О^ZQ�qb�t�!t��U����h�����d�k~,BUփU3�Eg;��k���g��9r��v&���E��-�( �����;Jo�R�	0�d[h��D�>6ѥ[�ч�w4�q��l�ߏ1��b��� .�]�x�p�u��ϓ�ʣԾ�8�񞪶�����e��:�f�>.w����0�D��Y&@���Gh���.G����e^����+�@c�|E!t(n�Db��]Q���u�_�4�mi��Hq���0b;X)΋-����Ar$~��f�D�\���=�r�WO֣T�
��V���V"7����D߼V��WB.רqV���g��l�h2N	s �{ 0f��D����Ē�ڏ�% ��rޭa�ml'�K�'�7&�R���7���m;C��.ޙ}�5_5�AMS	YC·-Q��9+��.k�N7�\���_��6��ܣ�Ic�v�A�e�&T�5Q�׌��5ϾR߲�蜰�5�{5�|��m��/�$�'��B�Z�?��f����gZ�E��>�+�m���~�=�~�=�:�Z6��JBͅG�ߞ��`2l��&�pxY�9�8��!��V���)"��q�9J�(%�#Obw�ud�^3g~����^n���(�e�ӻE!5lΗ5�A�3P�v�&�r���j-�$G��	�P�jR>O
�|t��E����]�R�E۞��$�:�����l�0��� o� �d�L+Y�I�E"��}Ejh�$�0J�y+J�d�M$Wn��{޺Ұ, ڮW�S
M�ݽ�*�4]�2��*���)��!�Ԉ+��K�`��ָ����x���6�nٖ��r��^)�2���{�Je�q z��:RZSj`vf.?9\���PyK�6t�-����.���Dڋ������lFFÚ���?�Qe�9c�qc���w��F��-�L%�l�~I���pg����aQ�d�r���'K��v f�169xÉ3���ħ�i��찰+~�½=�`��_.,�6��T��
�Y벜{s!�6<�k�B|a-g������U�c�,��<��?q<r����M<�W�[ˢ�N�/�8���M5޸���������k~���B��i=ز�(��b�͏�8��`ڥ����Vb1��>?����[81��|��g���9�N�`ϣK��0���/���Ñ8r�7loZ��E�	������K� �u���!�����@��t[���ލ�u&��$Qϙ���^��9�[p�r"&5��P�mg���Ȣ"�|���1�&+FC�5�;�q����i�=Ď� .v���`'� ���M�{B��6*Z4�꽱����aT�,?hF�3���b��{�yA����J��Yu�o���6��5�kQ�]<mБe�s������=v�+NS�>&��ڿ8:<ėq/�++��}�`k~a�Fd}tH��x	T<�_V��\���G�#�)���b�g01��G?xAy�o�α��}'�V�(j	Cs��OP1��,U$���>V +�U�����}��)�����f3�ھ�&=7JM�[KK�?���su���"�x��֜TT�ٌ�(],�}���1��c��n���W-�*W��5t浟�ك��~j��8͡D�Vư�A�>�>.�r��-��0���fsX�X��dQ�o`U��m�.����ag9�q�p�8�9z��n0�������W	�i��B~=��`~)w"gY�%���%m������y��8� K��w�V_���ť�8�Ԫ�0��k� �����O�-ȝES�Ҕx�����B	�`2�S��)�@5rQ�K���>%p��s즠	7u+XB�Ө]=:Na�_�D�kz��h(i�����&�������Ay��_��l�}x�'`d��EwTy�ecB�O��euz5huY<ķ2۲0�	���%�Yf��Î^t�10U@�����b@ ��y4��Y2�η6�aG��o���C��z|��o��/���>L	���/�<�JFmj�?W=��@�UCH�AnƝI��mWt��%�/Ү{��X�a�[#���3%Kd�]��a`�lu���!��&��f�7�*Fv����
F����z��q�sUcޤ��J_c
W fΛ��b�������^�lv럐.��e ��,
ϝ�t���c��0�
�䔨�L��CC��g�{1�21]���{�z�[��i���}@��*��U�o4r�2��e��;n�6� ~�%���܈�y��s���^�k�t@"s'���^�<H�����O�<Yu1����H�i�Z����m>Y�/
u�KuUlXUt�}��tj����tҩl���̃ތ`�W�?b-��Ӟ�æc�l�xU��A��il���K�I�3	~�JuP�| qB(ia$;��O}(J���h�&��}�{1o@����j@>�l-���`�x�r�{�:H�d��i�6k��ß)����l�`���w�2%�u����U�뀘�����ﴇ_��<�c$���g�|��P޲~�9�{ĉ�?6�խ�I����-�m�ـ�� @|����P��*�(ˢA�*���${���W��W8-��0B:$��F�"J�C��ARR�vi�_�U ���U/�x��u)}��O�Q0y�	�n�wo�zQA�/ j˻/:�p��<�q�Hs��r��xwt;�N��}�����^�KԒ,Q��z�h)�����}��U��`��	�bw�S�ʉb� �2;�^�߰ppT,�\�S�T�ވ?���RqN��\�X����q[*U��59A� ��(L�Ĺh�Λ�	A��! �P�.bI}6G��6G$�w9Z���o�����oݬ�߁��q+�,`�V�&۰�����
7�>��>��3��Ι�y:D�*6Η�N^�,��d7���/�d��jG�c����QҋL	Df�Jq͈6�h�.4~=����[e�0����Ɉ��S��=!w�鹔�ݺ�Y
�L����Z/�:�e5�0p�����'��w��ϙ�:�3�z*n�j��1���S�1�f$&HU%�!����i��Ό�J�k��t
գ0-jB7���75�'V�g�11����У�Y�r<�T�Kf�AJ�(hE�uu��@
l���σ������xU�ڞ����M�� 3��( ً�v���
�8,O2�1˔c�bG��Y���,]a�נ�+<ew%�E�Ca����x�������:H�*9���z |��\GQ2��/���섩�p�V�
\桱��ّ�Pt���� ���iI�b��P3���1-i0N�"Y�>�hap��ؕ�60�y�Gy��[+:��ݒ�ӳ ����Y=�h� c��.��
g"���}����\�d~��Ft#}�+Z�՟�� ��G �?���	���HH���"V�5� �!��qs9�ȶ�Y���}
���C�zVd���t�{=Ii7z�� 
���P�}�w��}�p���7"h�4eO���G�y�J3Z��]J�#C/o>>��wϦ���=.^p��21�v�n���!����k���#�tA���z�!*4bckF���ip���Ik��>��k�j��^!����͵�E��E���� ?ZOE"�?My�[���h�8Ǩ
�9痝����k��o�u2ﺙ�)�z�pO�F7����U<���.�D-�&Ok�/�:���~�$��:B�٨���0�^�ӷ�ZQ�	�lIlC��o�����iXp�y^��� ?&�x��H�(|2��N[���p\G9�eޅv<#8Y��>߄YI�҂�Qm�-��A��-k�B���kT�vGF���W��7 Oh����0͜�,��Ō�:���A��"{Je[ٯ��#��3�u*O 9���;4�F����3����-rx�*}�'��_8+&�@"��Cc�����^�Tԩ���L����5�By��/��5�C�!��q�]�ƺ̝��P���B�D� :�}I:`��F�4��Ł��۠��ғ"�l�$�u7,�UT�;��,̀uY���q�cDsz"�B����K�ߐ��0kSc!�u9�Q��