XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W��Z忸���`�ҷ��^`g��A2�t
�OSeC���0�D9Z4�nAb8ل��] ���2�c�-�uEh�|5�?a�N����i� �V��!�#��%��f�s$*�6��K������ߓ��mY'8����$1���&�焖U=�8u\�5
�_�;Y�[�*t!+�=�˄�\HTוּR`(/ze Gx��P,�y��Y`E�������w�}
Z��p�r�J��JE��}L?�Jg�٫�ÿ���S�Y7%ğ�k�1�;�7U�n]���PL��@�oZ�{ᛂK��Q����r�h�k���rU�Q�Qw�哀Xa�$y�V�B��|2��ԑ�pb��M�Q�<���C�p���K+Y�'>�\��� �;�Z���<Rd_���P�ǻ�\��Τ�����S�%�� f��èX1��%6�+q�$��hv	�����#5�H�jr����Ar�+A��8=�n��$\�I��v���kW��К�H��u7���X�h�%$��8sv��ʡ����o��rV��=�۔Y(ʃ��ꒁD����QhB7��۪������C|�Ճ��Z���	,/F��s~�Xm,-a����NL	c&��cT�ޤ�Aa�	���S�oQ�,����r���������хk�t	��g�T[����J �`�*##�q�@�㴢\ׄs0�K��go9!ʺ��6 ;��
�4ĺ�ֈ���X��à���]Ȍw� �u���bä) XlxVHYEB    2bb9     ad0V{ٰ�����oq�]��ak�$��8�����w�{K��-b��
I�<�d��*F�٦���[����G�bfr[,9{���ǻJq�U���~��T�����v@�ͫ����*MI<]ޘ��j@�0r��Td�곈����U@�?��Ơ���kK�Z�֩����)�2�,�^��ZBl�S ��z��z8��=�(�q[0��c�n߻���p����&��r� ��`Ց���ؙ׍*��#����m��4\P)��M�Jx8	�S 裷�����)��1ni�3�#��'9����h��y���#<8UYλO�8.�%3[yz&n��|NZ�Ŷ@�]<]w�7��}���ChU�5k��y���CLS�N9X�3R��ږ��og��K}b��0���1���V�_Z>9�[��|��(C˿��~iM|�r�P����}W"�^�U� D��O/vi��5�q��f�zĐu�\��g7��H�h���G�[�\G�uƏcQ}v�x"���0cM��"���M�Ο�1X���-�'�"�qg�!
zm��2��d�a�hD��?��_��ڡ�J��z�(�*춨 .`�M)5̺D�i�ؿO�}�T�@�%3��C s�r���Sq���Aw��`�������PY���\�K�p��Y@�U���VᘗO� �mq��,���؃���p|H�v/y�J���@�Z�%Qm�"#P!�+���]�pB+����úh���b�Ss�T6�imy�Y���nFl��ŀ���B��j�i\G�yÓ�.,p��7�+�J�Ww����F���f-7�	��j����@��璢�ӎ�*�{��X�k��*a]d�?��5/����L���	����FQ����C$|� ,;�~�t=󯛂@7+^�g���.���Γx��Mz2�\�t�n�38�&��F·hI���w�5G��sZ�S5��	]�7!�k!�Iŗ7k�k��V��r��8�=����/�UOW�y���dI-sY�o� ��0����KdTe�V���~ɔ�as^N�9���[�4���Qb<���z"��P�wl/-iCpC1�ކ�*Ë���z4ب|�UIC��B � �
Z$3��w�9i�i�{^i>�C},���gfZ�TgmG�^��7C&nn�Z�S�:�t�ݗM������O�H��Z��g>�(i8U=��Ƿ��'�M	��� ii �4�z+�d�u.��sښI���<l��m�9�E67��ܵ���R6�'�WpO�b���J�C�d��dSM�Q}j*����`�$�O) gF����/�KxY�|f�ʲ�Y��*p�!ΤJ�^��������[J�M�=e\-.4vl*$Zs�L�G`�ׅ�}��E�B��#{��
��#���!�[�� ��c�e�H��ՠJ����0����f�t�^�8�����e���t��3f�bG���S ���M�rr���O7h>��钣va{ERva�����f�<_(��\s������f���P}�O5Č��ߢ��B�d0b�ř��i�l��tٓ��k�;*}�-�Y~�gG+��9���_0)oy�%�����j�0Y2/���~ga��bäY��'�~�G�@rR�x3��,�����Z���-�*�ѽ4��D�w�����r��c���虒��"�ېsb�"-��+_5Yza�%��x��1u�cFJ舺"����-��WC9���E�h۰�qHү���Ȋ�GvWvN"S�͸vVV��TH�p���W�m��������_-�Ϧ���/	ݒ�6p6���xJ{�8WC�cނ�1�S�X7�]��h�)�7ş�s�@M�V�c����N	�˧�k�F��ehf�K��b�|�'����`�"ʋe}i���#��:����d��5M'�qw�M���GXçM�m0�H�~�Ӏ���e��zӘ'12�=���z/L��qM����`����v�����	�"RF��#�j氐�G�h梶�o0p��}K�� Z+,��4i��hc�Q��Ym�����4�g�ż?���X`�WP�[6z�/��rR�Ĥr�i�ʂ�*M�`��U�7��W �r(���f��Ƀ�u��k����Ƹ����݂�c����;&��]EG�M�K��y-�n��<���;K�29d(�z��҅�y?����-;����G
�:�n���7�s,�_�`�/JnuVY�۲$�J��;K��	4pX���|D+����B�p��̧ �Z�qJ�����ֵ i�����"� I�G�Bi�<��Y˼!�,�d觀��:;t���B�43����{R���6g���9@�%W: ΃�2:p�^ae�\��`}zܮ*�AZ)\�� �IpQ�aȘ�W�A�X�����F�`9!|G��M�=1����D����b��1���S\�ʈD�>��#�#�G�XW]'�'��U3~�G���=�1�j��6�ԁ��ǎ�Y5�������!�/�6o�!V��hd��%:`穡�{a=B)旕��Rd��®	S	12#�W���B�Fx��?�s�>~42jhF`��G������>�@�
[(�[&��0i��d֡�B��\����ɿ(�:��r�����\�K.��y�e�Պ&�^��t����i
R<�G�x�����%"(~�4ǚO!�O�MQ[-���&���o���`ض��}_��}�53��#lu+