XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����S�^m�b^��Ԟ��E��8�R��[7�w\���2a<���C�!��P��r��>��6����g3!�/�Z�M]T�y3�	�Q���5�A��'�%�.�\��iw)����פ��,�r�{�~8�D$Դiڮn9����ZkN�����_���r�;��rCn�A8O+���m��/���^r�7��+�M�c�l�8`�5�Z�S6�����}DiGF�� �X��N��6�߾+�5#���I���6���M�|�n5�y� o��{I��O}⥉ii��/�h���fn,-@�$f_�E�\]�i�Eiݍw������Z�8��gZ"�%Rd�I���e9�P�+z�/ܫvv�]�:r�yʾԀR��s/��4k��jFݱZ��Ṥ߲��,�cV
������7:l(��1M�Y	h��:���Y�Ra0�6�OJ�)�t�(��#0r��z��=�YT�S�9�&[���]-���������{�WXͲ��z].B���R��8������A��hDp{$�3-���Y���cᾌ�g�D�X*aQb�;�d�2Xt^:�1���!�P�Si��G�-h��⎓�X�t�kK��6n�K����/�c���26Hy��o�*�/^��7�7&Aj?��0�F�b�E'���;�o�X�L2F�zZ)v�Ob�Wx��e���ئO{X-�	j��Dr��ߎ͘Єܔ2�6�D=_�[�݁FŐX	.�����/*u��&i��I�1{5mq�uvXlxVHYEB    fa00    2d70̖I��Bڮ��m�� &�fn,L��`���(FY��wa��8|��R�(7X�3���Fj�)���6j�+o�G� �щs1�'���PQޒ2�8K(�A�����Z\"`�HmT�� �P����iY$W;���h��/-T�R$x��E��<f��𧻓h�8��v�J��1�ֳ�3M8��:��������R��rV^�al������)<f���*�m��H�j<�+Z��������غ[��USAc�Fl��9�
�k�̖-��q\	J�,�#�-yV�H6�q-�.bl=�b�������.�N�4��o �
{��4TF�J��^�8r�k/�`!��@�T��nF7�`g��d\>�4�LV���~�s�9BN������[�Ǻv�M���4�lifmD��J�5�2�}� 3�9�w���}j<`��XٳC<o��L�Ŋ��k�2�pA�rQ��;g[�:Ru��t��>c�E���Y�g�o��.��4��b��z��r�W4�~�ۑ���WXxU���~��K���%B9�����a�zy32�~/4s,�����ĬC|p/�U��RkM6��������<�0�g滷���/��1��d�$�j�nʨ��`]f�c��0���ҩ�|�td�wF�x�Ƣ`wcc-t�̓�`���˻�p�88��{6��n��-W�/��W
��0�C	��Q�j9\��z�m�!���ʇ��&��=�X�vO�/Xt?��.l��#X�/��{�8�Nθ��D�]��7�뫉&Ra�M�;3)�M�-̼+�ku1<S���	����契C�D|���@��Sq�.	N�t�nN o"��3e|��n��SQ��w�D�N��ͣ�͋wO���y�6aA[u�����3O��TB0��;Fӭ?C�x�>�Ν�v<�T�_$��������ߠ/Xy�d 5,�h��1�b'Z1����y�:��w~~���s�@���7�T��;E�Q!9q��ÁU��Nr߃ z;�_�#IwEY��|0tO��fjɒ��_�n��~���I�߈�FQ�5 �9�F��������~��#�e�^*��?8 ��$���>��2���f_c�C��	�~����H�LlJ+�悻`�_<~���7֐d�\����W�
�IV�!��41j{m� &l�	U���tV��9�X����v�y�IK�	fܘ���(�S�'�#��Ԗ� w4���Ц�ʩݍ�)(RHH��fL�ֺ�c&���)����^|)�5*�[(��QC,X? �Qu5ݻ7��v��F]f-in�� j�3-�]�v�O�r7p.&m{a��E�����\���|�;��(���i�cX�F#B�xd�+<�������ަ3
.!*P�~"/�N����JD>�GE��t�_�=H�R���تTc�뭴����s���(�� |��n�g9x1���Eވ.|�`|n����NS��FO]]�f����0�C��SN������~��.�{vR@g�ËKɫK����=}H�v�x�c([Rx���'�l�]	5��R��R!��3U�f�C�!p(nZ��������5]���c�n)n�*j�D|V>��~�y�$��w�,Y�2�c���a��ĐI���L,x�����ߛŃE�M�aB��|�� o�HpAٽM�OM��97*vg� "?�<���X0X0��4���\	`dW`8����э�f�HP:��Q�0VSt�Y��U�Y��>��jW;N���=�VU�9v�Yjm�d�Ў�" \
|^��ַ�Ie?�T$@�0e�?zlw�����e㗻�� �e����z�<d�-s�[gY6W*BM��������k�?��	~���j2�A�T�h7>��y���{\��!���JA��~H�՗�T�����S.��-�V��
�Ls��c��)!qi$��+!j]@���\\��?a\[��@m�r�/����}yj�E\�J�����9�|e�w�]���r�F�`�ex��~������ lt�d�=@��{e�<N�A��z�Ep����S
m��M�f5Vd�C�y_��C&f��
�:���we�@=������9iպߥu�ڻ����:ĞC�����R�S���ߢ�z�Wi8�Q�-Mr ��g0�&@j4�R!�<�+�H��9�U@��&���-}q���I��vz�جOf����߸�7	=T�v�gx��O�}OԤV{[���-65��UaW�M�_��N�u�v��Y���N����n�����l3�.ٖI���UAqZ���>�q�?��]�}�PO�D)a':Z��R�?�Z�8ֽJΰ�f�$��ܙ�_/~��>_v���a�8:I��|t��k"׊i��*�{��AW�EQ����s8I~��b@�ߗ�4�����aȡ4��d��ł	�G��̴WF0?��;���T�:K��	�:�����K�Hۥl�N�bd��54#T?ᶦ�$,L�F������Su��
B��F��	
��H1�.*�
���i����tH5���L�X��SA�V�b��N��&b�D�m���>��j�u$�����܊��*L��dэ�l@���</�H�kI���x�\0��Q��3׊2�:d?��\%aP� �G��,�v��<ѓ�h!��gw6��(=�V-����˒�Ɩ}y���t�:Q_�q��+g��ҭ��Jz����� �)�u %�+?�zɩJ�@��k�����:�������Pg�^ׄ���
?0С7�ȊnV�m^*`��e���:7-cg������]#�ZL���H(^-r&������>�uS���ӌ����(_�#^hP��t:Hq�!K!��W���V����A�ʍ�x���E4/���sڮTⴕ=y[��^�KS2����60:�om�u�W�
���2����XZw���ͫ�%�QR��AU��8��J]V�S6���fg�y�r#��N�g c���͛t��
���`���Ig,�O��q�������y@J�7g����R_��*�NkJ���.7�<�ڿ�����n�x�f�����}��0g�ɅC����9����5pH�%i~��N4�g�����Q��?�$�������J�Q����87��x.�0 �1b����+7�[-Չ�.8�Ԃ�ړ2\L(,H����ǎ��!�=��r?������yʴ�Qb7%��zb B����ئ΅�[����~���/�������a�l[vo���Y��j���~�&��ya4ʦ�r�纕��æ?Qp�?�^z�H�j�+b�6L�U���sLE�ȀS̆S�a�g�Y�:�," �Z L��q����/��s���^��]k��,#�)��;�lo�jVIG�5oS~p��{q�B�z�dL�\9��q^:����&1�|�8JD\yG��ɩ�`���-Zp���י�yեO!d�˒y4_�m.�S��:�ԃwu��]�<ќ�xJGD�,t�kD!<�vЗ�r�v1�GH>xvf��\�kHېmC�=��j�@�����C�v^;���q�<��_�V�ld0�}�f��S��s���]'�v�4�����q�m��m�0��`*�g~g��	"��������_���,	������('k"�x���W����p�fR��"��@�	�Z�}V\��I�X��4}�,�F�Oǭ*"*�����u���f��r���-h��N	yΡ50id_�Qa����@c����N�z�<�K=#����$�h;;��N�G�02t�`�G�V`��n�4^�o��ʑ��)o�U�Vu�
��Q�t ���r��y�ks��g�7�����҃λo���E_Q��Y�q�ˬɋ HK��W���dD��R$�!��"�F���<T
����>d��I�H�����������aV��?�� b�r#'̻e�
�@��ڗ�D�}���%YPt鱑�`�q���k�����ϵw�A�";q,�A�p,�7�C=m ͑$�c��N�����r\nS��0�n ;���ȵ[М֒�#�����z@1@�W�L��/I�۩��e�<
�Y�~��Ingd;S�h�Z;-��U&ϩ�ߖ䬕���Y�V@��9h�=�t�\iXp��A]���§�{�X��n����������w��s��-�U��1+��aݳjy�~�i�B�(�$�@`vӳU��G�:��>=pi?�Zy�{�_���b���/4��ӚY(�,�b�I�Ѐ�����9UH�4,d=L�<LR/zX�Ĳ����rH����v���Z46gvH��y,֣�T:�C�qo��
!�WG��8Q�:�w�*C�k�"�aW�*ӭWR'��MTg�{m�jz�QZs��o8'V�Q����Ǯ��hy��:m5�0�j�!܃��Z�1qP��\�+(Z�w���k=7Aa��
gғ�H��%�he���@}��
?�D����Ad���m&,�n���+���T�߰�@T��F~\$כf�CF?m�(�%Jw�x̢��xַ�W�����0@�=���H~$��8�1!D!�7�k�J��Rxd�B�*|�:�"埱*��%/V�S��N�0��/��P�����ا����K�9
�8$�;Gd����l~��	k��-��s�"x��d�GJB8��j1�W�΅YE	��*�ZMQ]wf���2�nb�H,��5[&zR�)qg����-�iB�W���t%-f�:��G�\�нg����5�8����zl��e�	�)�f��=hJ���?1��7r �2��טz���W�2.ps}�������nJ]���'�pɊFHú���N�ǲ(	~!��U��_¡䌊�v��ѭ��E_����8?��`	�\�>4a����;|��EST1�����E5"[RI��K�P�ޢ�+��*m�����EF�<6@�'YR�Q�ߺÕ\������7�ҷ\-뉉Zyg�D�XpZU���Q��)���
"V:B�c��޶57��y��aN.Y{�L�k�]��}=eQ즍�8�,qh>����Q������$zK����z���i�����kvE�/j�}gL5��t>y�����2rO� <��L��f�� �y���DbX��ޮ!��dj�` ��?VP�bZK�啹I��D����,�Vh�v�,��%��Y�.��dJ�ÍL����2ט�~Ĺ�c�n[ڜ�+(�-2獃8���C��¹%Ě��y(��ݗa����Nݮ�b��#�9zU%L`TҺ0�n�K����'����t�8&���)�n^��Nv��{R`�L��Ã��e��f~�>�Pr��t��F���CǉŹ-X�%����w�45�evV3��c6>{0����2_f*c�w�F�8{X����~�۹o胤36k6aby`�iB����NMOVbZy�c��)p?<P=9hX� �0���!ZL8ۮ�M�_�]˿��:�U�p�r�YE���5'�!M{59MX�|VC4P�_"��N��$���q�^�*��'>��/���sm��D���V���dV����]�.��K��Kv��Q�\�
	xPE鿖@MH�����kw��`�	��A�%d�u��U5���u4O��x��iH��aH�Cn�I�q���-0��?f];�ơ�ߴ+:�a$}�'�6A��}k�����x����W�L"�iǆ�RT�꘾��q�;qD�_��w�*�J�{�^�p,��l!o9�?��D��=�7�pGe�k�MZbc�'����@��,)���k�Z�ő���^���k�/�������y�b�l����S�\��^�e��_jY�5B�Wr�ww_f��e�Bl�7���7d�X���QSL�6*w�J~<��&����4�5ۢmxO�{y)��,cJ~�x� TK)�D��?�\;rW/�K��b,E���/F�45;O���:;��j���r��*^�u����Ɏw�L�U�zT�]8����ֈ�@�U� �(�a����W�;�ޟW��Xy���cсUkx]",�.ȋO�T?b<ܲA-x�J����cb�d�a�AW$�����7��(Eu�7���{�p�߈X�ݝ�;ĭcu)�4;�HWb��r�`
����w �_|�A��8F5$�x�}ьқ�� �LѠ�
<�61��S(�����vC��O������U��%v�����ݯ'�d�?��c���;ɴ�BM�U�(ĒhAY�^)u��ڨ]?��;w
*�X��V���U��X��/��G�g�C/�!��K�T.A0 g�O�?�.>Vlk^`����Yy�H��k�W��!����m ���3�m8B�V�ȯ���v+yl���c�,����ݹ���z�9����v	��Ҳ�Nyx��������9-���=����}c]g�?�F��KE� nc�����9������ XIe'�a]��=�S�{%��]�0����x9$@ɐ���T��3�4��s��s��(>&��N����l����������G�j3�k��_����<V��`Y69���ر(�.j\nYFn�U�c��8��=�E?�)($�HO-(x�cq�~8E��I
S�\{U��~��(�,������^$#���r�%Βgz	���<��ĦP'qo�ƞ�5�·�mc-�/-r: ���o�̳[/��P��@u69���K����5�뾷|��h&z����<����bX�[�=�PX*�u0��[WIeD���z}���zg�E����$*uw�J]��_̑>`_�8��A01���q�BCj�	mQ���iD�%���D��G�DRߧʔ$5��Ju�NӉ��!M7<�	x@ VФv׼�=���������
�½|��`u����{���6�,���!�=��T�6�N���9T����τ�"�{]:��y =R� ЊH��y��0�[~�U'D�J��@Kb?w{}�Ũ��,��9�����i�֞f���ͺ� z:v����z�����_�3e�P>�,��
R��Pa;�t�~9S+(���z�L>��[��]�����bX�qų���p�ML��#��M����13�=´�����a���~rBmJ�V$b�F�n^q��ӫTG��q`�28g��i�?c�9�����>+�}��9�`~�u��tp}i0]���{}F��m�u1���<	E5 �ĳu�g؛t)�Q�$F՝C�/�
�j(r���l�jׄ�OՃ�G}��B�䳇#�y��|f����� `&U�mq6��	�o���?]Z;O���Ѫ~6��#�!�|���ꝱ�*�\�<�	�e�WA33���Ƚ"Ȫ��}ȅ�����]r�y�W�U����A!W�0R��KO"�`��ぇ���w:~�$&d�)L��ϥ8�
��#�i�@�y��f/ӫ�S������U�4
h/��פZ;-�"��+%56����u2�^�o�1s��.9�ǚ�>Q�������2��WK�_3OI������b�t�W�CPU�c� �]ӗ˗E��%�Q�+�Ҡ���7j��wd4�gCi�h;u���9:�Ҽ�F�����ȮUv��דZ��S��wZ�PQ�����XĳS�_|��Ϋ��Ǖ��yҙ�9��"�k��U�^�5K�Kp�����,ǂFP�}A^�Nv�;`�N:��{��w�3�8?��K�3rN,Z%,@0��>����m�����ސ\_D'�n�w��i,��>kIHi۸�i0�٥��A1W�_k��E�ž AL~V���~x��E�N�>�!rZ^r�ŕ,pp��u˥UT����;ڲj%`n2��~3��34��<l��d��;�S�&HPC�C��Fo8��c��k����ޕ��)��|F�џqM䦿?ܟ�Y	���)�F.m�{��0�Sq���T�����2�]��~\^�T�>|@?�#9A6e6����~'�5�grJ �ۤ¾L����
���=3���t!j��hn/��2^��Ý���f1�0[s�P�aP�Tj3�m4C��!��D]�}3�f -=�R�u�\Ll	W������5����u�s�~��ͦ�ǅ��7�h5��/?RX��u3����$�����$ܫ�aǼ��@�k7��������a+i��O�%6�x��CH�����n�p�@qr���8��7W_P���ڵ�j J�)�=n"1�X:pEԪ��<��(7S��Ѥ���l#�q���"�N�"�8@!�[N����Ԉ�N�  �	ȺM�2�!mC�����~��0c��{�B>]��Ca�U'}��ac��?�(��LV3"K�$���ӻ�l���7	=<��m�C����{؈����P���4�ν�U*�1}^^�xf���uS�4B>{ֲ����K�@�<�c����̵��s��:f�y~ɟ�9ۢ1��1��#���M�-�ae�!D���=�f�1��C���/ƋcV0����`B�y� �YL_�%�%#��~�����վ�P��ܸ�%�D3��J*F�9+�Ư�D���~+��+� jDe�q�:�����./���<ă�'i
�ʁ9�h�J���E8�7�p-g�t��
G۪Z�*��os�{�&{-�5+�Z��G����q��������[0��{���W^�Q&L@[n%�0��S9��'yĦ�j�)9��jP-���o/�2
:^��z�(x���!Ϻ��$<'L4��X]�!h-D���`K���v`�1�7G�n�-5� VV4ĸԉ'��b��c+��vnx'>�:c��/Q%~[�XW߮35���RS��_-'�P�O�\��Ј���vϜ#_���/�*G����tg�z(�q���>��V�o��y���J"h4��-�.lQ�;��ݕ�Ɩ?+�ɕ)��}��s+�V@x�_ء��D��i\S���7�d��Œ��쎶w	����� �B��-��)!��_���o�f��,�qo��-�X�	G�3;�w�>�C	_��ߧt��!�����Y���Ջ5���/g`KӪ���BFM�3@�	�����L.��m�L��Ϧ4,��Q�?�ڳ�w��~�����6
я]�~�WF��~��h<��"�d�C�^��N��`��l ЇS��ӄ��3�Vd���y�+k�W�U՟cJ~XH��b���/������0�}ĵ7�K<��V?������Bw��}�s����e��̉<�Y��-�G���3�C��|u���8M$�m9l�5av=�6v(�Kpl�)��3*9g�uqX,�<{���y�$�k�"��^�y�*:��5gĔ��e��i���L�(�m��S���;�Иv*~����W�6�Mv���*�|Yh@�wG�}i�YYO"���R��*mT�
vm�¡O�M�&Hv�L�g��82̲z�������a�����چ�Wx�t�LMS�X
I���cSPw��$y�w�:H-D�
�p���������(w�Æ��d���xI�a��,gٿg�I[d�3jU�IL��L�Dʹ�T�G�L�R�6�I�0�ֽQ6���;�-��:o�Qα"��&�NqN�bHYy�t��
���\R�iH�f�2x-��`�y���L�+H���{1���r���=�c`��q��Q�9�{�A1I�g@������x�EjcI��	³�_'zY��S�{��i��?���ᕒd�t5�g�������na�ٵ����򆨡颤e��;i�TG�~���(#�,Y��?U�=1�-��0�)����9!ZѦ��c�w�U�9��������~G|�2W0�1mRa����`s�u3A>\��P��<vp�į����F�˩���;%.�r�g+K�� |�B��{�+O��ub5�7$�{ʛSa~��ԭsT��k�T��H���v�{� K�,��Q�� RxTn-�P���12���nԕ��f��O3�(�-z!�+آ����z���E����(��`��k�u��M� K\���揠�G��r�^V�0��E��ڌ�9��2� M9NL��5��?2��>Ӵ���jX������C�KƸ��NZ�E�=`�"��"S囮V1�$/KjO��ʟC�ud���.�.F-�Lt��H��b#o��Î\��^��W�Jo�_}	[\p�\��Cr��6����R��p��Xgz��pO8)�5;eϖ]TDh�=0GV����u|�t�_U�e���t��ԅf�DH]�&���P���������?��E԰����OU]IVfP�� %��|v�������H�\�X'�K�U���X���j���q�A����f[v�X�������<��b�����d)�x��?��-C�Y���8�K�J/%E,�t����4X�@p2�e��\�դ������[�;�[��:%�~�N794�x
7*]AiT�@h�5����`��O݄���F_�nH(�%������c�ڱ�m��5 ���d8E�ܶ��÷.����S5���TW�^[�dd	HR��c�\���y�Q���F�P�`��U^k�Y,:d���6����1݂+��C; �v,��ڳ]@���j,D���� �t*��w:� 3�ķ�.���7���/���q�ľ(��O�,���m��v�������솓P>���[�;.�j3ؑ�q@y���O���D��>>t�d])�ǸGf��y+d�!�5�~���	�mLf�J76�n5?ت��f��5>�B���tG�uP�s�̨�r�Ή�8�:CN���&�!�mqH_�	j`ՐL	�8AdŢ�E
V��͵�����	����:�⢛!Gm�bj˨Κ`�:�"�)�
��ڮ�/����6I�$�<�a����N.Q���oq�o��Fag
Ҍ���V�������f�X?f����d�HT/�Tb'Pt�.*������7�i��������qEr^���b�vD��k蕚O����P ��v��Z�[|���k.%?�uOL&��@ �@ �"x�V.CA�N��}�o�1Fm_\��U���m�'뼜ɦ y��`ax��w���:�;��r麅�.h=���+��K' ���=��_X��e����� "٤�_�B���U'�X���
wL*Ie)j�%W��"����>��<��>�c��Ž�*�?� M���GW��yq��Q��X���Vo��2;�No�WFD%v�Y$��[���8lu���� �*���i�s|��h�@ɝ��F� �jP��6 �i��|;�h)Q��|D�2���7%���<��Ć���*弛J�LLv9� (I=L�C�w��rt6]��?ؙ"g�l7𣍴!��uE���d�@�ߋɰ -����퓞������c�,M��c�x^�o5���"
��#e��i��7[�����"�J)-I/t�8ϓ*(�.��[�G!Μ�XlxVHYEB    5902     f20;Ij\V�ԩ�ȷ�D�{9��j�(�tGr���^ʫ��0�a_���,���@��z�oӇV�ʎt��/#��^�8�͓@<��F�p_�s�
�}�� ��+ M�7�Z���)֊�.�[�[#z|+I)��+�H�:�R[Q�
'p����:���H��5L-����+��)�����5?ɀ�#�2�v����ǫ�m�Z6M"@�`BJ�F����Z��V����һ`�ա�:s�S�P�"/�J �l[8�Q��DJ����U���#>�"���c�M�-�2dV�M*b^���0�{�S����5dF���Rk�[>H��_|����P��bP�9����C�\5[cL`b<T	��V�Y�Ut��lrߖw��x� �;�Q�6s��mn*�ݧx��N�K�B�>�Jdu�����P��6pW�{|%U2�:Ao�'�x~��0��,�Z۬=���k�>M�*�y-����scCݭYԥ��P��h;BR�/�$?�����2�[+���O@�O
���G�A���g�9���5��#�����US����dM��Q�ܣs�(����J���E�*!����g�cP�*�&�OM�����$bv_k�|r^��ϑ���/N���?C�~�iɌ����2�|OX�\�;|�����^���\*��R�r��H���><�8�0� �'�sDs��9��2��6����S �Vܦ�o龄���/eԄ�*yּ�@;���2J�T�Q^�b[��f׭�RK^�mڜ�X���/]#TF7�A�̰$?���4 ʶ<��RX�������%��\��~ǁ����x��)*��
e���[H�f�1>���������P0߅�dJ���7��2Nؗ7_�8�:��$o �U�"��jh):�6�Ӵ�k�㎓A��1rWӥ���:�
���Ɍ���X��������^nU�.��,�����	48��933��4��1�2�Rw��/�ȫ��r :EKb�;�e�Wͧ^��_�gD���ڶ�v��Ȍ�O����2��C�'��kFl�2�<�(^��k>�`2��G>)�ٝ���/S�lr,���E6�ؼ)��w1Z�z���*~�w�֮�H}i���"�y>�zS��~�+�jM���k���'�E/z���p�>���cH���n��~���"^۟��=]1I/Q�P��f��q�Q�������Q]��]ìz2RT1�#�~�%�kя�������;bcj���4p2�y��cc#{�bbEZ֟��(F�%,Wf �u5�*�Ь�F�1*��"����6�gb�l�������RG�@��?�l��s�JM}%y��"�3�v�	U?b���b|�f}��]J
�4�8q�kx�� �VۓS�=?�K�U�L�����b?��|�e�աi��={Z�G�Zo���F���m:]4��Ŧk`�����v�9��~��Y0k���9��ݕ����w�����S��P`ʟdu~~$!5V;j���B���g1e��a�U��!�w٧b��x�f�1����i�nPfǣn�>��ʄ�z�v����9ζo�V���
�BA�X��_���J�%����������n+�I�5��s��F&2�8�z�ek�*z�3/��0���EX(��%�m�r�����f�XF����A��Ԣ=��#h�ʦ�epA�9¸fY����ܜn��B�I������X����"[�QJ*�Ym)��Gq��ڠ��y�%�7�Q_.�<�������p���V�:�R^���n�ą�0%=����W�&�tQ�{������L܃�%�jA>rݾ>��d�(���]�ɻ�?b�M�)T�����eR�7푘-�x�v�g� 9�R_S�J	����>�Q0��J}��L�v� �è#��rd$cu{9��9�u�H���{�^����̤��n��!]�I��|�7�av{ʨ��@C���#źԭ����41��y4
�a�*4��L�ظ�~Zr��f.(��:)�U;zPx�:�!V+�@���*�F��t��UҾ� 
NX*v>��̂�ɨ��x�<t�w�lD���Y�����	��J�FK�%+�r��#�j}�[�EF��.�l�% �S=�Ӛ5
��;����i�*iS�OМ=��v;3%�Ȼߛd�����B�߀AK��6�1u�Ԩbx��]��TG�KO�!�h��N@p��U(�y������*��� ��vp0���]X������q�d�((�z��yZ��;�q����>�ӳ���y"/�,gɝ(S�t�K�^�xo�o)	ԫ'D+y�u�tN�X��F�^�Юu�n��>�q��y�I�\�C�n�:��3p�F�E0�������..�	9��6x3�q\M� ����1�y��OK�6�Q���.�>�6P:�N���ߗ�*�6�˃��$����U��B|o�;	�V���A}��W�&�VM��څ����%3�b3�������=�U˫���4:l�3���\�@F�G���4]��m�)�Z����5����a�MM�nfu�xe��W61+c��0�R��G�t��Pΰ^~��]n�s�r� �9�{R��W�BT΃������n��I�l�i�(__���ɇ�ָ��g��+h)Є(��²�>2#�|p7P��cN�%Lq&�u/�fϪ��W��~LA�_CU�5���X+1ڻ���!�t ̓W�r�o�.�B|GH���d���<��3S;	p4���n��^���v��C���>����C�� ��q�'ُ8j�� �˰�B��S��=A��7���]ˌ�g8$HbՃ-u\�+�m��n���}^߮�>F�Q)���Õ ����]ъ��Rcw�G�:��6�7��A+��F�(UC�Ö
0��%���5Ep��5��V��Ti��9���-)h�b�tO�߈�y<�&�2��;����n��6�M2�г�Z�v�\(���z�
��~�n�:�����,P���'���'f8l�)�*PV�OW�o!�X��HοnҴ[�y�;r�]x�lR8�
����bNI�����B��^<���9�[~�ra�i�p�̓��>�w��r����G��阗�W�ߌ��-Uh9�4������l��?f��u�	���`���_ ��w�V8�g:�	;�E4��t�I�Ä٫0|�+3�n�Y�EȮ�����r�mшb�.��(V)�o'E�O��g����l��N�klP�"��OS�ɝ���u�������O��]h����6���
[D�$�r_�2��0�Į�=6KK�#
:��"a��СD�e��WP��0��11�!�^Ӂo���_����џ��5�}6MߜU�鋒D���}��>���W�!�5��Z<h���a�o������l��#�oE�ދ�z�f�!(s�5����U ž���5���m�G&H��3rνjƯfJ��	�ݩ�+�a|�|���6*He��7M���^��(�{�4�,9��T���)��+un��)��0��v���|o�j��LcV��[����뙾$�?���r8��ŉ%G@�!a��M��TJ2]�F�����3���$����D�9W6���q�i������L�~�n��#R(B��y��(�P��ns�@�<���m�rg-G�Ȋ|nr'�J�E�Bv�E����BE)�i HVw�I�"�B$Y��l��� $�O[����-	�Go��ոDw4^�g5ǲ�L�,As��ZN%���z<�($Sޢ�f����G!�賞�������ՈEV1�ڔN��ر�wj�8�J���?n