XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8N��!E�(Ѯ�^�D���ΐQ(�B����q�p5f���d�	��q�=�K����E��2��E��+۵}F�л�q��=(>,��=�i����T�#�2qtS~����P�(6�I��ր-�����WY:��+���,�}:���M2�&˧�������
��[�U#<�m�0����;bY�r�����4e�ު^+����ts����{����b�7��g�044�#W8w�8w��q�]Pے����B;�8>������Y�ձ�w�
�-d��G�5��^Z���:���ŁJK�yL�V���[���2�r`�$:�ը@;�o��{����e̤�$��d 󂑏�¤��7��X�Ib�ܠTdW_8��(p��ڀs��Gz-@.SV�.���2l�����X�9\q���(�e@a,�2i^��Y�r�q��Z���`k��4`*OF)�m�f 9
Yv�'���&k 7͞ܹ�4S��rڽ��u�=��Q�	���#	���!<L����V4��j[�������a�O0?�.�� 9�4(�U9.B��_{�#�0��,�'�Sw������s4�)�$��D�32-��H��2�ض�s�J��`09W��~V�#m!��܇��n��S�����O���f�̋�s���QQ���5�ޔ6�y{���c�6�5�<4&M{%�a���ԎA�Ϥ�G��!9�7���b���÷��{�-�v�nZϝ�fx>�4tO�Buj�Toޭ��Z(8XlxVHYEB    5cad     f00%��R���n�e��	.Y,+�ĆS�y�i�S6�~T��lW�&�q�CKI|��7�v�S~�xd�5&���T�p�Rj�^����r�����3Zr�z����1������h��>:���&���l�=�pyv#�qK�+t��.1�~��jԣ^x��������άF����칭��3�R�֊-C�s�(�wµ�|�D\RώuM| �H�f�Tx�ӫ�$Nϟt�zỵ�vH����٥ߗ��Z���ܙ0x�;��(6&�v�&��QC+�P�`:�0Be]�O�d��J�%�l� �k�+&k�+�XاH�r��P�#-�Yf���!�`����O2��mq�m�9�b�����^��P�>>`��������g_�	y�����$W��nE�2�e�y����RYX6��8-����h��+����(J����Ǻ�\e)�#�<G�q�z�Oo;ߍ$@I��)ÙMEd/y�����vD�$G�Ӆ
�Lck�ⷥ�
^� =���-S�?���Vaa�#���Q|/�J�uk���(�k���v^n�h�1���>��6D6��!V��J?-�k*��v�U!��ŧ�MT(<Ԡ�E����;�H��X���s���Di���!f9�⇎�Za?�h����S���;Y2] `����~]G����K&�j<k�	؊^��lx��B�0q�$�؟��� f�������cO�G���@1�B�ʁ/�Q�5\s�^�����.�虦֋ף@�m S�w�O�
������_~�ys�!���pT�gb��[o��K�,�x��|5|�y~�?�R�}*pU�v-�W�+� ������%��W�d���%�����^��_��ʴc"���� ���lԧ�n�y�.��l(X�*H |��2��oؿ��c�A�D�%�L�vT����`^|��h})��ү8B�jߏ�W��� r�<"��˿q+?l��Nau�G�:��D{��^��e��|$�P�f=����9����P �=^!�C]���*��d�ب�B���|X�����_���ͱ<��9���+t8QU������(	�ʨ<��v�v{��8�,���l�?B�����Z%g��t q�gE�s�g/�g�h��JV��5�eA_���G=_�	�,���Dm�������ü��Ɔ��3#N��k��j�̿J6껽�u9�6U
w�\��r�!�c��䏅W��o�q@�#]7���f�k.Py���Ƴ�D�m��#9[L�@���`Y� �Rw�#?��Y�d?1cY-3��(5�X=�ʡ~�)�q�si�Bi���A�}z��9�F?�0k��Xr��DɐH���8�؈<�
LQ'J�`���xh�����j��ƥ4����}�1��j��g�dn��i�zp���6�L�_]N�U�n.t��荚"�-�8��pM&ʱp/ޕ�H�M�;�����*_�2y�͡rC�0�w��}���lH�w`�QB��dq��w�J��x��� �B��5��;YP�짂���6^�	���m�و�%�SI��/���|�
����l�Iګ����mϫ��,��qQ�i���+�a��E�V28�V�x"�L���{`��g��qA
��A�9�]��1�=���_ݪ�ǻPa�dC��!�e'"�mv4�����F���E��`F6i���d?��ű�
�o�GO�^Ha�u:�;vZ߂dQT���k��H��`N�	-, A����:���%c��`:t�!+��5FoR�^�J�6�-o�طCWO1
]=��p=�d_rٳ��<����2�˫!�RB�|N�H^1jz���x�J��K3�f:��$X`P;���f�� ���iӏ?d&*f]�ʱ�����k�ڏv�m���(�m"Kjx�s��Ƈ�b��>Ѫ�A�q���$�L%o�M�O?�^Z������/�\��`
��Ϣh[�
{�"B�������r�H�$>E�h�E7NݱH��:#Ii!	���Ms�KPO�3]�hN�~y�M���0���'�ɻ����Z���wZ���q�
�_[�4�{����E8Be_7�1��׳�!��N��ތ���o�.6�7��VV}$ϻ��0?���x�dVW�'	����c�fT�S�h(�~�x���c�I�d��0�Ս�#��1q}��Ƙn���[�̫]Ua��߭�4 ��;Ms�i�VT�PMq�jB��$|6��L{�m�&��P���o�7H �U�9yE+��6��fM�A�.�h�)g۴�[(����\a��T��	JT[���^8X�&(�;�N���c<+����1۽�E�h��i���~�E��?��O���^�\�Y�a;	,j��M�i�y��,Q��W��ՠ6�Ӭ�H��2r�@��X�o΁�E5l�S��g��L��=���h$ �cm�p���l��괊�W�OH�?X�y�M~���&8�L��5�ŘJC��.N�Kͽ�ӍgI[{lE��4� )�֝���>���0�����[5�ܾ��r��P7" ��Ph 9_����N��U�I͏�o��
8����ҚW��;��I��=�z��0�ܓ�����{�C���oz�Jmhz^1�N�����t�j���V/A> ��~��v����HS���w�DK������-]��RX�L��=�cUY�)ӎ���;�}MTSt�A_3�gT{��o�$%v4E�@��Ξ^�
��{�����qX`�@Eb��3��^� �V���(>����E��Xp��C�<��Ag�O���5�Z9#�	!���"yo���!B��CU��>��~��_�yʹ=�f|�EA'L
*��c�yB���lM���b4�.�b6��a}��Gax�w��g�(�N\�(��x���w���SN2�P�c]�WY,��0��}�cj/�dϙp#ęM�bp:w��{.T$"�!�DEK%�Lu�S&�N�]i�E�L�fHԵ���ة�"�w��̨�� ;)�#8>��aU��s�j�"�-{�0Ʃ�M���(��߯z�����|s���_��Ր����)VT�8�����t�*'G�b%*�It����^Yc�-W���a�h�T��׉�X���ھ[���K�a�ˬRN��Ϋ���^�o$(q�'�pۤT�!�'-QJS(����x����i:�zT)�Aɲ�h�r
�*�vA�*�ݢڪ��=���7���	 ��Ⱦ�����}t�!b�-S{��qS\�Pz�Kq�dy��~谂���f#��׌5�a#w'�	�aE��tzLp"��0�,����!��<��ss�i//~0�Z� Y�nM���}L�j(���ZQ>�b��������$���y��E���u��Q[���W��Bngb�zF��/�����[��K��p1;�宭�*���3��$��^O�	q9VB�\tcE9�gj���	�96���[�2'b,�mɎPn�A���i?D����B��/��~�N��(�{-VIB��?G3��3%9���-�\�7�� Jy�\�d/ڋ�\L�!�~^��c��H���B^Ǥcּ���O� 6�8+�═�g
s�[�3ｅb�rI���#��cZi(/�ņ����"6����d�)o��(2��<6��_��(���q�I+��Շ28z��X�}J��x������o yS�w91�D���T����ȣ�r@H�ʣ�U�oNR
������<�����J�����A^=�N(��Gww�rp���Lj���i�����:�su�H�l�p����