XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j��fٻg=���Pen�䝘���h���x�i��Gw!�� 3��W�"�Ü�VM���Ȝ� ��|n��-	��	%�Ǧ>���tj����@"`,>����6�p:>��Ϋ���Ѭ��.l0@��B�c\8R@A4���W��m����p���=.ȱJS�������$�	Xߺ���j}(��A���h;I���g�\t�T���œ�����Dagli���.Ҿ�k��7d��[���@�*QB,�N����$�5�s_2=�N/̔%�:@x�ݫn+i�e�l�{q|��޵��I����G*��aZ!h �Kw�dq�܌1���g� ��Q�a�ΩĠ1y[�<��O��l��ҧ�ШF��� ���09�=�
���G�� h��(�w���� ��ė��#�O�D�<��O�I�x��:L��X޳[���H����bUK��� 
gq:�����$j̺������2.�<oCM5�Bo�.$��������w��E��A��#Y��wR���D��$	�4�
���Z�m�o���kl���m=
���t�h�9��zp�-X���C"�}�vF�c�"r�h���$];{o��vx�,7��J8@�&�Ԝq��Ѭ��a��Z���M�3�Ɍ���ٝ%����$!�4���^�X��MN�Td�_a�����|\�Y�,
�����)�cR��<g넳QCƬ����L�����A�s�}���}����3�3�h�XlxVHYEB    47d1     e90��ދo]�7/�*?�ƻ�1��5M�֜7f���d[j/�ƥ�����}O�t9���"tם��c��rh^�Z�'u$����`�:��"wr�J��k����C�Q}F�=،���X�-���	���-]x��u��q����x!����S6dK��3���d�F�!|�p�9�/b��Un������P��陾Qjh����KP^1<���ԇ���Y��'�Q��(�tV�P[ܣ�ğiW�Xz������W_\Nh��j���e�Jk�5�ސ�d�6�L{k����Q����ͽ�X�5�(��ߘ�䃔n@�5J5���kL���!q���)9cU��l�����������V�Wp�p"kۖ�|�M[Ҹ����Q��
�q�$I<�,�	6�Ly��*�fje�~�a��Lo?kf�ӿ��y��[�6����ʮ���M_k��)#J%�*��F�߇��K�Z��a��*���9�z��Qc��N ��{�ηq$1g�%I#37�*#$�ٸ1�U&Q��)-Gb/���,���U���,�WJ>���A�Ra��x�xSMJI���o��d�ϫ�4'���"��j�$�%;P�Z-1�{� ����[�J ��o�/��8�[�jOM�7��aN��o�a뭵(Z^�/	�����,g��d㓶�O/��f�k�[EBW1�M����!3����z�x�8��!%�ӂP{��ɵM��e3m}�g-�&�߻�A�x�����U3)�lU2d�4#-	�(�������"zv����� �w>vdVִ��ć/~����?QP�P&tk;��6�Ih����{O�/�ʼ��3e $��	�kَ�d�3"hJ�dt4�I�q�-<�1oT��s�O��+d��3Ғ�J��y����רo�+�Ѵ�8l\����TWG@�*��j�U&��TM���Dv�:m|Ա�!�x��G�Ǹ[��G�$GJXe�t��gA�a���t�w�5��6P�}S{ϊ�B���(״+l��i�Y�6)6�8��6w���Rb(ʸZt�~S��rd��2%pT��a����n�.��H����BGr���TX�͸tī�|�{��ۜ\�萑8x^����Lx�v�y��< ����W�:B� ��y͚F��y:uk����I�z/���/�zSM����v� ��j������ʓUjU��6����W�	��;��1�|�g�CH(sf;����4t]	&���a(��;�<J��w��:8�{s��c�	T��د3O>~��4	Z� ��r�S��p
����R��i���c4XQ��x=��1���N�[j��u7����\W;"��bm�;�\�����(_o!#xM�-���cq��W�����}n�]B{�81? ��K��r��:�!RC�'ퟥ�n��WؒQ�
�QJS���%����9��Pԏ@cv�Ykr킥�T��<�V����.����yr�ϋ���Q�O����X�X���H'�����}Id��� �$ձ��zA
�<��9�h�r��l�z~9����J�;� ��`�X|�Ru��mS[T��p�Ƅ]����%����5�r�$�uM�0#�ų�ϒó������6�ʸ����
N��J�vG>?��덕��`Ãf���i��uQ*�B���hI u��k��Թ����o����cƻ@D�|�\?��[��sՋ�.�̥si���e�c�[ھ��	RE��I;w����1���C�^��Ҕ[�:�'ne�o���le9P�H��B�[���L������e�p����5��4�SQ�}:�o��MB9I1�-�-�ɖ>U��n��ڵ0SI�#�03��FT�*�����(�>{���<E��,:��T�5���zb�Ĩ��e��xa�:p��y��u������z8ғ$BR��}�l���Jd\9{X0����1�'�ِ&1A����	���|�yƥ~��K��?}�_߶Jd�{���cT�x!�5^�M#��� �uH�N�4Ag.���KOL�AbT%�t�5�)훔���tO�ςfȔ�T�xU�s�KR%%���k�����_�0�z�>�Y��vji'�Z\�bp3�GC�e)�n�/3�4�]�Âƙdg��+������+�;|��_�Oh/���awx�j�ΞULA:�7�����Wo�_�<�@��b$�}�\T?�UE�rs���ُ�8ʫf�K����.ǡ��>M�SDCK���x{d(����ď��_k�n�2ğ}&&>y�� �8ߎ���q��#E%��ut��R�Z	���.���
 ���m��H#&*`>ҡ&[��M��9�`��{zd����h0��F��'u $08�2�������Y���^(�����L�Z�u/�Ǉ@��ܜ0鄌((Ԉ�ۀO,����/�����,�����K)E�z7(ϋ$�W�}�T�Y�q�k_[4�l��2K�vd��������Rx���ݭ����N�����k��r|I�C7-�~�Mx!��6�R�Q����
D�-`�r��n7�U�T�ה�L��<qG��*#{ʀr\!�>��&��	���Vf㜣���:$�q�
�>�*��9"�8�[��~���ިI�����.����	�1�Aj?��WW%���]�i�Z�*��ŗ���-x|����)y�>���À�cj���y3/�^������l��eE"fRZ2�e�Α�V�ص�|Q|�
T���C3�h��{sю��D ��쓽�֞�) �`7m�pD��~G����y����r�.���?H��������D�����@'�U`�~��$7CJ��ÕC����o� ��9=� Q0#�����AN��!/Ho�eW��V8���&"�ft����k$��2Ԝ�Bd,�Д��t���L��̻��*O�I[�,�X?���
'xɁ�{�v���`��7�(|H��^{5���$������}`��$z��řC�RDB��ž��W�IR,v$>�������V�(�y�$�7i&��>z���ɂ;�Q#���+�JJ��c���:m�$n8;H4ο�c>�C��X�<��<�_Ч0d�\�DZ�G����cbm����)�&���YK1�R�g(sJ�Hz��aĸK��K����6�烋#~Or��'^�K�Jj����`�ú����z9�"R�~wY*}"�
\!cĪ��;1GJ���=���J���D��1G�*M;'�_t���W.�x(�쳻5BXg����������tO�>{��;��][y�1`G��?�>Ճ�t��M� �YI����M#zZţ>�����0�,j�1��1��H�R醏=ui.��!B��ߒ��wd��=;x9I���Ŧ{��4���N�;����Px�Kf�yř:&*���&�_���5���ôs@J���SW��|!C�6�`����/c
���e̢U����F���տD��1��TC����E'(0q,W\���ٟ��h
�(�Dg�����yp�P�Zu�V<�L��E�"�X�r2��m[pH[l�mJ�-�b���G�ޔSWҗj_��������T��@��^�6b�QpզY~�u<y�}�5���Qϟ!����q��D�f-E�,��

>�R�&�O0�z[�Ad��سG��Ef0��