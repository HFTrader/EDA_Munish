XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/0MCq��s'?���Fl���{��Cfc4i%}�|��kt��;J��{T��G�՝�]uk�� ����D��6�A���2��
�K�����On�cn�a�ѠM����	�u(=�� �4�1��~]����0�0M9�&]�t���`8;Z�ITUx���9Zf;ܔ��^VUbnfI{�Uɩ-�������V4�G:X���C�'�=:����#�	Oǭ�s�|x��޲r����OWƯ}/!Ж�7?;���"�LF^\Z�,��0��{�&�Jߤ�^+���(�p"f0tj_�Hh1Fy��˥��@G���z�P�"�����NS^F�3/ �En�g^,/��2��-~��!��ZL�A�IaAN�r{\�V̈��M
�Y��?�^�9�yK��c~jRZ�ri2yp�L�x�_�B�������!�A��͚�
��^d��<=H��Zv�Wz�x.���nm;��[���OV��M�R�-1h�-1�A�'����@|��(QA��e�1'�#w���8�.��l;C�W7/z-({�*-x�ę��*#��N��5���C'�3U�;���#����I���;KI`�%:Yhت-w����#= P
|u�BqQWC�e�Ji¹{�!Q\FE۠���wp%�Qm� t���4��/gKB�?Y�
my) �&@=��U�B�����"�75�Je(�D�5�,o̕;���"J��mi��Ƙ�U���N�n�d�{v9�`5�m>]�Yv�Ưa��p��~2��XlxVHYEB    42ae    1110#���h6�g+#���=�I��$o���Ü�41SACǺp_�{�5��/��pG��h5x+�U�����`}��zۆ�����2 @�`�ҽ,ڻ � � (ClR �gx��ɖeO��^L��-�\Bg��(݀�GA��6�Q����=Q�DM��X�]H�eC��\4�ێ��ǀ"�t?i.�g�5�*0C<�{ ����Gke��J�
y��zZn��)�$�v5S�B���za�Ih<��K�d�-:/�A�7�k�yC��ୟuh_|���[`q)m�25�/�i	V����
�2'Rv�ǐ��jF��^��S�U�cW�Yܮ����z�L4ۿ��k���g}7�a����jr�!�O��%�> ����)4y���X��;!BY  ��{js!��0�i�I*�*����ةN�b}1�����z�`JwM{����|�JĈ+�P�U8>���^TQ����Y��VF� �#n�����1�D�,�*5��U�����X�sV�zXv|G��kB;������z�����r������1j�쳴I��`���h���PҢ�"�Σ.�x���*��a��ݭ~)J�f�gCZ�:Z-�l+l�(����T�Z׮I�hL�T���/��g��Q��ct;���Rcq+��&��lrK���6�Lt���\�y���h�A*GD�	WeR� Fw}"ЭYU %�£��,�����)�z�D_��ح;��e��
�#`�w�2��� _�{�� iҢ�;��,nK�2i���^�-��?��J���� k~ƣ	�2U6H�����~�)#(�4
��妆P,�6G��s���r?�R��yO����(�#)��u�W糎����\��X�����.��j��E�5͆0SC�f�9L�B�/�������\I ��Z4<3LPۂ�y!�4�B*n_��E�Gc�fk��o9ü�zd^�t;�r�<)�tj�⾿��>��-u�Ec���v�-�1�I]4K�\�^��OW���tH��m+�[���~��_A~���}k]�M>X���`��b��/�č�),�Y�c^b��X�LxԤ�`�DѺ|\���ۂ��EU9 ��?2��|�1����FK�`\��m�|�0���=e�/|#S�~8�;ɾcң`������1
8�T�Kj�D�Ѫ!D�}(fo���:���U��Cm����S�ǒ��t�`x�w#��7�57Ʈ]�Q��Ba�������Y"��+o�kGCB�n��9;����!CS�2rFlY�$�YƁ����N5�{ ��$K�a�sYr	�{���h�y���v`jI�Iv���t�J�߭�Uy\�w�6>yo�(�������UQ[|�A����-���|�JH�U�=)G�Jg���J�t�Xq1u' e!�}�c�+U�k�N�m��́��ê�z$q/>��(�!D�з���N]�܎Θ>Z��z@Y?�X�jI��������8Z8V�S^&h5�κ��h���&���3������A���x�D�W��]�7S�/(b�a�`7�>uzP��
�"�F�(�s\O��(l7���>E��80[�?�
��T�����J�y��/hÎ虥�f�5��B��گ���;�I��c�5��9� �`�M�	�f&-2��J0�4�J�O�\Q	$�6b��ą��U(�l!�ʬ��[�~Y����7~<��H|�(���i	�-����HI�Fta-H��N .tu����v�Fn��d�1m����[!j�۹��p������P�J\��_9��|����n�A��WĀY�ts����j�h7�¨B�m��QO"�O��݉;+$v���}hQ/b�XﯷB�qo����u�*��}Ygǧ�u�J��n ��F�R�
x{ۭi��5���D�'��I�ΟFo̷}U{|-I"Z�)��^��s��ND���[��r�jX�4�Fs�uվ���dz��o��:�&�(Iv��1�av��� �,a@��ۚ	��$�2�WOyR���=>*����ps{��{����bk��U"͖fw��7/�(|{Ab�!Ͷ�*	�=�����5�P�m*����	��]#�Us:��S�%�N��jM᤻�(�b�4��M�,
���/�B������)�V��8��mf���5���;�4֘������6��卜_4�`�ܼ`ۓgڐ���;9� �U��c@�K�V�c:%r�E��*�T.�D�p�]��Ѐ[���$��ŧ?f
O���Inɖ�k�V�)�,��X�����8c�
1�z�ׅ���!��G�T��.�u�V��w4^��.���yHZu7RCg�f���Zu�a�#+� ��#�]-*�3��'�O����?������YtOE�� �����d����x�.�u��ҢmjI�@�;�����l��U��w�.���>5�Y�/Z�h�~��<,K.�,�wg���dTS���P܅��{�"S#��x��2B�-��� ��{�U���(�x��PB#��/ns&�P�#�%d��c��� �i��f�U�e�~�,��G0��z7�� <�:`aZ�$�+�KH_d[&>�!ا-6�c���/u7��\y(5G�l��Y,)vڹ�B�����7�Ow,��X���m�	���̤Wޤ��$�����@,�@S?���h?N����X��0��v_���?�T}r���+g(3�v$ך���'�K2W|�U��@�Z��Cf��2)3�^���K�:uv��i���޿�}��A�-��$�˞
�_���� �1�e�$�{B��/RȐBgh���qt�O-BD��((_Eϝ��ɘ��4hb }�B 0�����n�
��ph�E8��l����P��A��p%m�8%�	��N�r���~P���Ǵk6��ߎ�yd]x��x��Sy��Ģ��O�:ސ��"_�I��{Q5\\���߱��vU���p;i
�rAB�I��O-�m����#�E���1���F��4�CM�]�$��R�'y]��H+-�V�>�P�+�t�:BKVL�d}��K���_n��G��1�?��/@?�a?v���Q6Y�zF݂r4�r�#$�>��Z9�qe �qB�������:��Ar�R}���#�WsS�D��<�=P�F;����#��H�8�[ʏ���O�@6d���:�Mw�~�1�}���D8Q��2��m*σ�U��%Zf�x3R�z��A�o���N�r�����"�u�`�@�%Q1I��r����mM��� �뎽����3]D��v����'�����?��� U `��7�����Ɂ�Bc�W�Ec?��%�n����s�g"��#��@�4-"鮦���3������*��P��o�1��t�s�ŕ��64�lj �@��P_"�1�ȠP�g�T:�ٻa --�ԳY� �8�d�������	i�bj��[�:4�S�<{6SY�7����#	O��xX�V�8�����#GL��C	^q���ל��h��L��f��	."{-��w�n�i�Bh�y�$�n�i�=��i1}��0�%ȣ�*h͂��#���g&_���\e�ae�bV�D�m.���>���3h�^̀F�)d���8��l�n��.<��R��Қf��Q��^�ԥ�̉�w\��b�E��_��p-.��8����h/o�|�\>zyVD�K�����	~YG�P��	8�!��c\��3�)*9�'�]O�K��i#6O���u�j��@��
(g0:P�x�g�o��.;_�m��ÒWE;�z`�����پ��h�M̰�+��~&�vڿ���ξ����фUXSο� �9��E��P*�%@�D��z_+�! ��-[�櫓V��0[��й� ~AUZ�� t"R:�Y�{�tO�A(��v��LE���T�ee��ɦ¼��B���轲D9�7�[���H&��Y�WL_�0M�Ltc���i�b�S�1�zwI�Í</���f0]V/����?7�v��*��H���8�7)�/�Y:B*ʶ��I�s����;H�7�?U�~2~M��W:O���{,�D���G]�d���u��<�����a�ׁ�G	�ɽ� �d��n�f�2�2� �\Hm�'���ݙhs��$[<þ�)�����f�l�x4���Q] ���s�Ρ��h��W9�j��v$%��d�&��]ѓ���d��gz��\T����ײhq��_r|�\{67'��]��maۅa5�B��:��ԡ\�����-�aJ�h6^��=]�)�d�