XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����[l�my.x�	�K���1N:�ۆKz�
���(r�o6{Ni��W��na�hNS�?0@�n��@�9��~�G��~hr;�@�����E�i��z'�!<���@m���&"�5Dm�㿽׼�L%��@�ӱ�M�O:i��$JZ�/�x�&T
�D3������p_�EK	5/��ۤ�I=�u���#q��]Rn�� e��V$��c�Q�t��ь��Z��g該͋Lc��*kQ}��	!&^aj�e���	Y��}��c�R����O��w�
i� ��\���0������(���]n�n���+��X-��Y�@��d��Wƺ�mZ�����erlDjL��u�G޸ ��c��Q=��E^L������^�edՀ>��r��� E����k����8J��ycV,���H1�n��ne2�E&��~@$R��tY��u�WA�%���|l�SK,���/.S
w3.U4����w�G�s۟�$K������X*9lYt���7}8$��Y��3��jC!��{o�q�m'����EG�}�j^$�d����m|��0��
z��Kgֿ	}�h%V���`x��͚2�4������Ș�	V��@:��M��,�F#a��Z)0�u���G�Ô���s\D�ؓ��^� ��씟V�wʵ�Y�"�Qm�Ҩ%^<��r��9��L��G�Ի60�+��jV^�4�6�@nj�~��oŜ&�TbT�i��Z���9<��ϧM�9���ap0f�]�@(�&ُ�v���0'�XlxVHYEB    fa00    2480X�A��$��ʕ��$��
n�j�{���j�g��iy j;�ܦ�W%�'�cJX��/-xې�oDT�@���"�:3����m�	����7���Y��uA=*l޶���w�K�0;HEQM0�/���i���ґ3V���D��ʈ�9p��q�܎7��^
��@K5&l8�&R���=A^��Ųi���Ơ�����	t�'��sU���TA���3kF���;G��Viڇ�x�j- ���[�t�����][��c�YuX�[xW��[�����M����E���'{��xqQ��0I�K�o'�Xx,�4��;��o�AgLƮ����
�˒�D<�M71��>c�V��ře�3�k�^د�\ɮ�#��h�-~�~�N�^��90o���0��K���'7�{�3U�ѣl�2�ozQ�sa�_۳~{��A4,nSs��pQi#WL������6M y��&���&Rv$J�W��
L`7���d�Q[d�̃�=0/s\�ۅB��ɢ(�(c�����8_����=�-��m7>�ι��{������_si��C�C��!.�ɹ�ě]O,��a��l^;Sq��(�*�e�W�����/�MN>�ܮ x`� �Y��Ƹ �޲Op���~�tx�X����VȄ��^a���R�%-��<�c��VLӃt|����t)G_�-���Ncguн E[$ =�v�y��f̮�L�6��x�
Pćo/�t����8�9��ܦ��� W�x�`�Z��t)^��+4W����o�	z�4��G�k{`֒�U�&�amb���r[�볔�g|��K<#6�y'�J��P}2Y���X��{�*�u޵�?95�k'n��{�PGԳ��<��H� ʒn�[����P�o7�ŔFf&��~6\dD�������8=�-�ա��0#���d�{���c���a�D8���ʞ-�+�R�^�.��C�7����)�)�Z~}�eR�cj�ϮwƎ���_Y��RG���U�1U�O��`�ep���J������N������F<�%��䢱�麞��DSspt��h��V���(-��t��������}��}'�C+ȴ��� �wѷ05Z���G*�s�&^�-H]Xh	]*������$B��\ڠs��nt�ee���9ѩaC�>zdM���1��b�N4�͇�y|E��p�ՎH	۬4[�Q��rz~���*u�
XR<��{��q0���LV�+�邦n6�������ݞ����]�b6��!/� �D {��lRI�"�NK���.�4g苁8�΃2QZ��a���� g�7r�gj���]��2-3���a�W��j�K�r7P��&��E����0���A&�D�3[�~�jOo���n2�D��S� ����x�b��]Z����A�
�g��p�3�����Z6���[U`��B���]_x��|�:]�:�O�-�C.�9�Y�m[@n��"K`���/�d��k��L���(/z���@?�O�&���c9�e�7g~�t�J�u����l���J(l�ŸZ��>���>�)kO����&p����7�
�L�#9v�ԔZ�P����}}Y*U�[��1�7unu����hTRY�]�+�2"7'R���rM��\��"PdV���{��6Gڍ/+�rZYee�ć��Ӳ@�JL�$o�d�Z�]�a�I��Mqg$�����X~����-�N9�m �_���������b=�����F@(�ϋl��{�v2���rg �d�L��n'M�]�8�]��<]�5Ȕ�V�yoU�;ʞ�Ei�j7*4�V� �@�nK1rmw�m෸�7.�`�ޯ�@R{�m�K ������,~<�n�ļ�ުBrLd�JzZ�+X�Y��jd�����]^�rm�ժ��zLc����b&d���57�ol����'��?�������:t�\�챳΍����mbp6�
~>���<�c�0���f��
*rpa�� ��{�Ɵ�g�`w[Cٳ����N#(�/x�૽!`�F/�n,�V���K�M[(f/�HfΡ�'v�JI��>Va�:%�ᶁ��y�	#8��N��.�w�M�.��3�r�^a�*8�`���=�At_�ս�J�m6��U�z�+P�'���`yћ��bѺ�a��C����E��6NItm�`(K�t���9-���^��@k����Yᴒ��m���n��i�7c��z'���$�"����ОJ��Tm���#j����>MFē�o�
���e.
)�W�f�4N��e|(Xt��,�ֺ;&�2��Ńɺ�R��/�Qcs���&�x�|�i��i��ii\0�܄���b1��f�_r�#V�Y��U8��UX4���evE��D�������g�@�a��pr8+O�m�rX�(,ɰ�pBP������HϤsM�v݌ڛy�L�p�F%z���q��ޑ$��������AG��d�� �)�f]�iEx޾^{EW*��iu�u9��rB_�$�+\��e����isǥ+�^a�*3<5��KlڡV�ߨ�Gp�8h&�;'+�QR�$��Ulw{Y����_�o���"%���M%k&� s�x_((���K��O�I͞Z���N�fA��4�1�9�JvQ��f	#��p��D'�f�3Yjk���^E�`�x�%��Nѱ6ļ���I��ω�~A��L3h�PvӇ=�-�=����2�I�s�+s�\8V�������3*�'����Du� �ay�@u�34���׍6d�C�OB�(7y�h�Xw��������S�c	�-�]계���J��J�Ů��'��D����Uj˔9����ĝ�*�,�9������с�%TQ�}t�Q^O0�/Ck�!E#00By��E�y��|�-��X�+N�k]ի��O�����?:������ƿ�y�Q��W�=�b6��ε��խX��9�1T���R�x��04����`"�5.�T��8H�i?�	䒔 �x[_����}�
 ���{ב����i3��t þ�z��<:�]�&�H�X�������u���2�Ҡ4����*]㺼TPqm%�ueh��KL�N��:#v��=��(��W�-XhvQ�C��xS�4X�ҽ���Ht�U3������E�ܭ���v�(�7/��nWʹԥ^zg��N��x�a-O%�S�z
�jDz��O�
�j]b�Q����E&�j��$PKGa�|N/��������c�{� ��7b��/��(T�s�B�S�H�M*�4#�.�P���
?[_�/Nk�2����|�#˶��a��T�uT�C�=p��r�5U�ʌ��S�����:U��4�ߕ�NGGq�Q��� ^R���!�kk#�����F
�c|�q��k �DmQ-�!"�SF��k���L�2��1R���Q�ߕZ�����:�UfHdU��]�Dg˭��^5~�A��}u�D�z	f���׹�%"�t��q��M����K��f��9X�)�#�F�k�Q�[��j�ψ�oJ���ⳋ��^b"�t�f��3�̰BV�gXc��^�m4��
�H�y)/*���Gdb����J�����X�V}��0W�X��p�ߐeV3s�<>�Y�I�UE�]/u��ڀ���ۉ
��p�#W�Y殌���.Y��w�@IG2o7���Q
`������N����g�H:�U�R}ō��:��!|��`���lx-^=�SE=+�R1h<�Y�cy}8�C�(�pᾟ;��YJֶ���>��F��g��UF���g�����MUM'0\��K�;�ü�F�qr�{�t�j����20^��լ\AA��/i�S� ���湃��3�#���
�Y�S? Ԅ~QmZe�I�mD�̌r�H4�+�o�N?;�t�`9��������/�q�U����%����Q�f�U��󝅒�����n~�з"&Si���Y��n����bC#�\�zaG�%!����g7g)"���'9��F8Q1*>φ�ȱ��O���[�pE�1�&2Dg`�+�%�fQ��uΪb}��x��X�CWC�Vb��5Kv��T.��mK�`�F�F5~� ������6w�o���9�9f�(�������мV�.��td����cq
Yw������:K7�H�[��H5&ȫ`u�_:�o��EC/u8M�"[ W�DU<���@�)6�`�l:�i���B�z ��t��j{�v(�F���!�q�1�8)�[z)�<?�JcQS����oO`��tR^���������uC�}���>A��;�R�ko��hͬ�^p��� $5��(�$���6��o�ڕu[�M˘��#.���0���]���hr�J	���#��KG�@�������4���2����7%/ua�p�0xv�9�v��D�3�"d�s_D)�	'b���ڊ��F�.��r������+���8+}�I�%:W�`���|r�wQ���ksaj=���؊�5r��>3�Жݨ�l��9�@���R��RG!v(m?�݆7)}�=�P�i��vV	ki��a��H�!�Sz������yG��=���PӺ|�0`�4�`&�u����*��M*eG"����ŕ��ؤ���K����f?Y�4�h�s��x8��7�����պ/�O����"[K?>8���2�Z�*����%��E/	Lz1�H���A����Z�W�瓩��v���Ed��gDq�aLVSLO�vn�?-��g���$��R��q��I4�N<���� M2��T��X�;��l_O�7�a���q�K�����UcK߳4 ��������|���@/t:�2���dh;w��L�W:����%�K��=�~R�!v�֯�[M�+��)�8M�)���e�J""�S��1E�����!L겶،�S���:��l���W�2q8r�0�����G�F���u;�FCڞ\zs�2��.頮*���[����� ��A~��%ŝcj���Q-��1���)��Y�ѽ�%��O ��[�:��>�1��n[yz�np�oh��?���ۑ��F�ښ\tM�*���c��|����X�w1D�J���L�+��CI?6R'�a�\�)|6�����2z�"�*?զ2y��o*��.�X�4�/ytG��CSP�C�:XMF�t�_���\�h����v�,_c�qH��n]qG���_+VU���2��ȧ�5x��SمN��|�L��O��)��!�/ޕ����4eG��a~(󣷊�m2VoIy�G�߾��[�C�P7N>�h����I�`�i���g�����f�tU .M�mX۪c�?��V���П'��^��1�?e#�����0�1����o���я��V��.�r��嘅`g_���y��������ٰ63�wR�  @H�cUKJY��m�Ӑ��0�9�/y�`�TsB=O��in����v)��OrFJ]� �:����\>=�Nsw�;:Fb�2`(z���������ZE�3�֕�!�\����a,��_ʬ�v�i��ۈ�N!8G6�왱#L��L�:�S]m�XD'
����A)�E�d��R@���@%�����i�� ��ކ������?��{��Z�����9�ڑ���!����K6o1��$)��osx���W�'0zZdY_�XSʝ1�X���,¨x#��:v�:�T�p) <���G\���"HbE1��zi�=άnJ� (N�;���u���:���DO=��)�\�ͳ�g��d�c�A��쑧G��]ȣ�'��`u��F`Z3��4שT HQ՚�cޛ��\��D{98!2Ќ��4-Ol6L����%����õ�d:r���� ��W��*PY��[o�ym ͜5[�>�D�$�3��<]L��e�_���U�շ�۸|���[�Es��!]5(���C~�=����=�r2K&��%��G�~7F8�w�昔�qzO���%�b�s��Re?s���X�ѧ���bփ��`$��W|x;������ ��i1;�Z�~�+-$D�Ytq�/IbI �g��f�鸝����s�(DP�әB6�9+�
g����stl���V��u��7�-�<�G��o��l��wX&S�+Ь�J��f�^[�W�*�\���M�n�Sf�7/�
C}q��1�`�#������R���(�������T�t������6�1p�F��X�F�gaYI��K&�&�� �Fo[Q�e�f�`�	=oo�2Q~w7QȂ�N�\���p�޺����Z	.(IO��)�/L���*A3r:VWzR}Zg�2|���<o�{-ƃ�v���u�C�V���a�a����)����~>�CO���G��)e���RސAʛ�e3�mp�9{���R��<�J�^c2\���o�x-i�)�w%�޺IWg'o�K�ڥx�T�Qɼ'��`|��4��	2Dg����g��*G֩�+k4�6�DKI1*�O^��)��FFC ��9��K"O��-�.�Y�b��[��Ϸ�-fZ4@�6�"uÖx��k9hea�f�dtͨ�X�ׯ5��/Uqj��'뫗�04֧1�8��TQ��>.�UI�J/c�AI�`����&M܇E�[�˛�
Y��N��l�3�J���c�ip�����e�s�(����8ƇڄI
Z�uӗ��-f5��4���k�AR�K���Q��a�ʍ��1zg0uk[�ÉޡZ)�K��~:4]����6t�ť�������^��K���t%H��{Zʸ�h�D�l}���3���&�Y -!B�A��;(�ٌ r��EӜ��L��UZ0Ҩ��:�z�/T�k�B��#�a{����������R9ӠO6��wջ��P
�H��0�b�=�����1u�'Q;>��7x�ܠEbu�?��KI��^{��E' ��WJe�,S�H'���TU���1_��6>^�&�/�r2'4H͒�`�m�����/{�j+�G��W�Q��`��I��H�,���wz�qP�4��M�M�n�Aw�X�.@���nZҹϻW;Y��8cX���٫%�d�u�s�l�?�u;*��' "���g6^[_
��uC +��R�|ғ�蚵��rw(Ԗ
�՞�Q���0��!�@a7�[���V//9d��g:��v��=�q�U��؅]64�J[��N+�8DZ=�X�P\��8��QE���$���P�Ya���Q[�K��8���-���ڀK�� Qn��ߌ���V	�Ukb�1� �z�+��󋔼#�M�4��ۡ,�����=2"z��
�_���&�,�4]��w�����B^�7�e�Fc$6H����X~M�d�)ؠL��;iN�Hb�D��4��^�-.�R��M�;s�v�[[��(�w�$h��-+|-�}*DK�G+�� �yl	��_)�ߗ�����#ɸ� }8��u���9����IP���|�\�"8��b�8G���4�P�,�%��ǩ�U ��g#o�}�lx.cG�yL�o��{������͠Z���̂1��?Jk�9��o����Ki2�j3�A��D!])���{���o��T6��.��W
�&G8��|��'[�]`��M���-��c7�&��[S4uB�'q]+�f���X�2�L��[�I��w�2�H2�kؖw�	�G>�<ug�7@��,���Nc�G�ǋC�c-Χ�D����*��V��B��7v0����
��r����;���CĻ�[���t����VT����kA~����	�E��JVu�1�"�ౌ��qH�H�<%��`ȉ�����N���v�Կt*X
Od_v�h+v�=�L��T��֠��
jPp`��5�w�S�<g�7>1!�����Ǧ��������O���������\�#2��xa�Mi�=]}������n�5$DL��R��3b=���f��������<�v>���8�v|�M~�4�W�T �.����ަ62��>�<>*��47�����4ǻbfh���5$�9Q��A�]�rW�(�i�G���Q�H����� �ei-N�W�R���E�����ػ�}��K���1kV]G��޳����g=�}@l�C��j�m%�vJ�h������I-l% ܜ_�z��^@�Ǭ� E���.hB��Ju]D������ĭp�U�[]^�	�[�c)�G��훾\]V�`E��p[#���9]�r9հxG"��_����E�._S�/ ��(�%L�$F
0 ��i�PA5������[J�[���&UzZ"5�I��h�B���v�d.��0m����"4��am���>�Q���J���a�ؗ���%-*��1q����Y�׊O�6*�K[{�y��)��n��Tېh��5~��l�Ve��H�/�3v�c�i��_B@���������.ȍc��sO�)��-���c^��m�+��`W+�8x�sq DKWN�Z߳MJ�n�~8�XS(S�kFx?Y��B.�[(C7,�w!���h��� �Y�Io)��ΝsT��?+�9k��.�*>�]�6��U�O<�橿�-5t���k��@j�)4�w�x3�YI#mOڦ�9ǈ���B����S�Zs�
�@*x��v��	����bΉh��__��}�UN$s#}8g(V{/�3	�K�1����="�W1�H,�c�_|zŢo�
 �H�rxHc���)��V�u��H	��ľ�*.����h�#�8�3�����H��s��!p�NMZ4�u��$9�f�fR�3�M�~�����W��4z�Ս]�Ef�)���=K��duʂ6<�:S���)�<"Z��7��
Ro�!~�����>d����<�rF���, �@m-�Cq��ĩ@��*��yt�2�����-BI݇�BU������Ҍ�tNU�"Ģ'�rד������)���� t��@���ڼڙ2.M��dשq-%�3y��VXQx�8��z�� w���}�
2����8���՞���'����3�r���n�|(���\-���w�����r<S�x)OK0O,1��[��7sG��&�Ό�O�C#5xu��ڛQ߬`-Gn�S�T>�f�8Y%�f��!#ր�%R����O�}َn��{s�҉Yh�=�+���%�H
Y�{��Dl5�K�D}���4R.�.�G���w��74��f�'9ʄ�A����
+�S�XlxVHYEB    964e    1150d!ҝ�0 ����k��1�|�y`b�&{����\�\IG4������rؼ�y|%�?��Z��X����q��D��{������/n�_۝q�� ��5f��k�Wy/ �x۞J6~Ao!����>�����N�ШX�&�J�"�h��5èF����Z`�P��_��7��.���R���eݹZ����.�Y�΂=�� �SDW#�6_4,T�Up�թ�h�r���B&�����\�M�䚣���f���S����>�.�*�9�;�	n���z����X�U'q���O�'բ#od��.ӹ���\�A�-s牄۫o��(�B�����0U����kOm_�4�m7D���N�Vx����qW�*����E�4%����=�Lh�r�[���~��0���/+��3��6�V��炪����5��`W�j�XGb��x��:��}���"��2�=!��IM���eb7����I� ���#��H�֫��)s'�o��el����7<�'g8�Խ�!�2�Pk��"?o���Ζ`��b�t�P��͐vꦞt�V�ͫ/�W���q !���h��b�ׂ2�0?��Za���+��FH������˧;������{�n�׮�V8��Z#�L5I	l������@i�/OQr]1%�U���cև�a�5��LK*�n�q��
����E%������mn+��v�O{C�ÖVd��%��)wF^�E�5o2�+�?߶�#}Z*;��B�����($2�Ҽy�R��4�j�K�Aڏr#uvs2h9hbͭK�C`�@�M�53���V,UN]�s����وd�;^�$Cd�)�����m���@vwe�-_鑝ו�o�L}"Zh�H�2?�QL�l2�u�!!C��gߏNS/�U��5e�zH����n��q}�;��us��X���#�:�~	ۅ27J�(F��V���G<1"�G&��_H�D�sN�Q��!P�@A��S�S�y��[���郁�XL��)�3��[��,o&�y��N|Ts4�[���n�G���HrG���o����<��,k& �q�@�'�[�|@f�$�4&�%��z��p��YT�p6�aSh�{
�e�]t)J��w�wf�c���
%���=��+���nlfv��h)�K�a��vܯ���	�ă���{�	�J`�m#
�h@�f�V��N!?�[��6�(K���*W�R�DH�K�:ㅀ0�.�q!Ȼ���߯N��e��t䗦;��^f�l�g�H�Lt��|(��3�X��Ìq��i���k'�d��޹�N��jsĔ�!|��/�UA􂴜�Ҿ0�:�1�#X�-.������7��T��i�~c2%_RI��x��Ŀy�[�����)�K�W��R��N�	�<��c����2����s&n�)RJ�kk��M�/(w�'���%-�p���5z���N];d��*S�i=i�^��Lc�:θ�V�PJ�*}D�F��z)
%���a��yҷB�w!��@�܀��(��vm\rF��y�[H�('L�����kyL��A��A��@ږ������܊�vs�ĊZ��#b]��ņ:����A�J�H�P�B��l#��v
���aXܢ:���	"��cM/P9�wt��g��\�<�ٳ���@���7��5�G,��e�.���zu:��Ņ[\���4�U��ݲ��Χ�*CU�J�~cn�'�uq�^Mܾ �"�iD
�T�D�>�ZrJ��C���飢�l^N&�#�r�[�vY�w�+�VG��.+a�^�g�>^ ��SF�6:�?]�Z���5�F�,)����F�7� c׆nA����V	8�kc�|�_�bZ*o�u�Sh]�d֤���nN����:N� r1���n�|h^�y�㖈�H��'��(�3��[����!�����h	+��K�ۧ ��ك\�����7ܴ"1���Q-O�|Q�:�l#����$�8_�q�v��^�G�L>@E@Vi8àB�f�+zm8׻�4���Ū+�2�iR��N�8���#�6r �e����Y(�;
q�X���^Ί�pD��+S�P���$d{*M�����6f�<=��"A��RoͰ�.{���4�6/��H�`{M��:� P7?�t�L�� �W�z)��5��z�_���񞛴�JP�e)-��<㯮����o8�;�����e
i;{hŏ���?��l{������띜��2V��j �G؇){J���u.�f6�w����9��N����[����h�k9C5�㸄�V��+�`�hqH���J�V�
K�>)���r���\�����NsrJ�������0�C�8�쀸�ӄ���o2\�c�����&dR�b�h��3Ů,a����yָ���T�g@��r>ys.v��~@M����S����9�n{��0o���ÁOƀ�����>3|&��p�R����6
r/��9	P�W;�R9�����l����"u{�����:���n'� �WSHR�O(��LZ ����AG[����\ُ�׾u:ڗ`71���s8 �u�w����#����� �E8�O�9 �&A���o��O�#��T:G����I�w�E䭼����t�l˔m{ף(�����n�	�#�\|3u��d�$s5���5o/{�H�6I�v�+ò	�2�B����"2±��N���e��Q�ẉ"��}��1/�L���*4!j?ԟt��s��+sM1��5���O�z����,rN�����Ű�%o�ш�M�wQ���Ut��[Ǣ/�a�ͥl� <�L��d0�SX�$���Ctv��Dw�e�*ᰐ^^]�B��`�i�\�|����#�q����MO��2��1�;e��k/z?�T����bP*{F+�'M�A�@�ȋ��6�գᾆ����S�q�{<�v�y����X�E:"<�{�F-����ې�W �KF�r����OE	�bz��-��$'뛹g��2a�7V�6M�B7o�h0�&��u�X�-�I�����:n����c���H�\2y��m��y8�*�`d�s,<���ï
5�؀n��3o����g49X�!�| ���q�b��#�H�`M�O�k�f�
���Fwc�6�7/���$4�A�vL;%wF�v��Q@6{0�Ǫ�˦;	��9�Ks$�/_���oG+[��7�&+p��y�F^�U��TX%ЁC�?���EKZJ�f��1X���ZjH��fW���r:�%P
c�^��g�7=[�����T��^h4~�j�Xb�ޱec$�6��4�oژ�	���^�J����"ͪ�����)�}9*�i�2�ń�#��0'�����wR���ղ; �N�SX>��o����
�9��fy�J�I��%qW��D�8͸DT�G!���M�'�=� �	PZ�<k��=��!1���D��LA;�+C��B,��NyH�Ŭ	�5���m�$���[P|� r�X��5��  ��t=����rI�
,�"��o���b��(Q��@��^d2$�g��a�%t�o�kuk d,�h~C�#'/l�E��i!*�����0��<;ڌ1��{6�90�D���窨��"�X���8���.E��\Pi����Ӣ�T�[�1��h''̫X�%sT�2�����ȅ̳ηO�%���3���jз��ʮY�1p}Tq�a`���0ut.fIx�<]gs$v� E��^�dtѤ�9�M+����<-j��&
Z#�E�Ƞ���5SV�Z��Uc����0������ظ�6�����X$�$�mݐ@E˶�|j�3��%��s�8\����P��7�Ѧ�����D��6\T�5�$s��(�L�Ѯ��8�F��_�Q���-� ��~�rl�"����m-ڝ����A	P_�� �\��s�Fn�6'��LCDN��}���d�tњi��'�Ş��p'J���OGڮYq!͟�^��rH��5��\���
K[�Z���B�E�=Eko��K����i�3�arRT�Ά@��z>j_2�-��M�$צ���z��$��� ��b<.W��zi���<�e�g��]!��m��ͿD�Y�t0E���#6b��0~��;���z�%:qD��7u\��6��%a;��O��̋���ǯt��r��j�`rg�<"�T��/�S�-&P,�u+|{Q8���U�b��ې!ac��{bm�ժBQ�=?�s�5��;�]�ÝfȰ�(+�'�d$��]�4���>y/�ϛ�F��˺�1�t�B��!�(L���QaQ����0i���`r���ᨫ�'�~��a�{tL��JZ*U�}�V8X��C���>�(xzt���&�@�L�2�u	����rD����