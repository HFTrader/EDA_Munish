XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ve������0D  �֪�}Ϋި�$�\d�rH= v����џɔ5�^��Q�j�zc��<�<E����7��>��Ll����6�#�����U���A6TI#�eжFwòwN�B�(�g-��G�j�"��8h�G(v���j{�S2޴A����;,�'VH�d 4�>a�Jp������1N�]/��(+�z��� A,3mK�N"�4J)0 }Rߥ���E@�V*�}��-��%]�Cn�Þ�1�Fˋ��b绵�����ojO@�e:��A����4�6����	n�
Kg�#��R��������g��*_m���`���虾��ݽ��*R ⊠(8ށ��Ⱥ���}�99�A�C����P��O,H�[�W�z�[����o�<����d-M��&A�R�k8`��1�U�y$�T�����5L���=}�0a�Y�@����ߓ���-�~o��%`�kxp+�����X�\�	��{����e���j1E���X/���􌮝J7�Omሜ-�C���R���G�g�����D�; thuK��i�1�'c��u��Ic��|��/���6A��y�2�IM1��5p�U��M`��P+m��:���[N�ܵ�7g�[~��D C&��Я�6�x�fc���f�IS�b�5�-�
j3C���������i�I�go1&m�ϕF�'�������>��	�9�
uh!��'�uc��C%�z�V���3
c�@䴙XlxVHYEB    5073    1100*��V�]Od��$��Ϫa�P���Ȃg���,��CSm��?��Z8<����l���3X���L��^�?X��	�nx�+��ĝρd���UE��������66&�`����O��WT��l�r�i����x��a��v*kby�C���@�0�|�@����K�4�u�"Z��ĀW��Оbͣ���RMiO��L�&��G	����1��Gͷ�W�=̃���|����7o.|R�WV�����[Lpm��3_ש��c�
6�e�8
PӜ�X� ���W���p����m� *gu���12@�ݗ?9s��V-�W9�́�9U�a�n���vel
e�1�M�i�gg��a��^T歭�T�-�� ����:I�g�9�v{���\l�V�b���3F���U���&RW���}��ia���O&KF.P"���t/���뿗cU��C��� �����Zc_9	�2��r���(Ȯ,�a%��~�gowS�֋F�%��-��I�M�;���6�_1�vuH)�s-�3��׼8C��)�eC�ޠ���&��Jʉ�G�0�e ;6�_�E�d���uo_9���,"�qp�>T~�ٹ+�����9�{Rr-��x��-�|t�	�+�k�Zd�����_@�S���HW.���m���e1L	TK*���t���3�]4�t'kʧ15�8 ���۶o�a��j7ne����5�ɬB�^S#BAC['���E]�P\T�╰Jy*���c�>�"��_H�TYK�������g#�K�e���6"�)X���棑���k}�o_~h��4�^47)���_��$�G���m�,�8�c����Vps�}	V���:�>���d��ڿNd�D�a4?|�De�}�|{���٢P�o��sQ"E��$�n)�-������Qs1h+b��E���� �/v?d���Qx�r���[�a�f:M��UT3����C(ݒ]�vqy���Ż1Ŀf*�/�Ji*ߏ�NH����b�Q�tC�<�>�z'����_�G�&?:�>�yӇ.�76�=T=�RQ�����Z�A��D�e%�SF֎+͟�L�9��%!f�]�����Y���,y��� ~q�\�tWV��W�!��_�f��EG/dUb�]+A��8[Rk���v�Y��C�ף.����G)g�x[�aW34I�'0��P�Y�Ցb>�u���t��*K:߯�u@�����዗;ã��Z8��N��� ��ln��[���}+��ކ�,6G��Ajy�4:�G�<�� D1xj�0M?q�g��gJ �h�o��A���S��ཌ����J��_�G�P蚅���-��F;���c^_�i�\������wU���fL�%�/��)X���ռ��w��=_F|{���� ���S_R�H���Y�jqZ�F��4ޙh��,{Y2��"�lE������r�*���(x��C�in�E3h9-ۆ�g�,�$�|3~�g����������I���v'��,��x����~#�眦�D�ጩ�bAD���.����U�n5$��E��E�TM�־p���5�[!4�d�4ja1Q����}���Αsh,��ha�W���k`�؈Dz34�W2�d��t��5�����u&�]���?���+����%-�S\V��҄~�$�U��۟H�;�EIVY����r���U<� -�NG��9�Cp���Q_��ۏ�,WPq�̩U5a.m6��KbQ�.��u�`��y5۩1�	e�ȋ=:�QyI����7���AB4���� ���	���uT4��g�s����R�	�V����vO�N.�"�p[�6�<�\?=Z��7�>�U����BϚ�jBn���K�"DR��Qm��Y����^3F����(+[� ���W�W��2;�^�d��<�;*�WO/���RZhltB!�y��ˣ���N$�[���@�p�g��:)PmK�U��:���g�T�A� ����9g3�V���-p~�F=�^�]a�;�o�oz6
{*������X�R�h��YDQ���)�]D�8��@�P7ea����~��������:�l��}�+S&����o#��I]��2)ͮU绒K�nh��~4�R��r���A�u�P~��G�1I�Q�2� �Z%������z�^P�Q�(�#�Q��i�
s�mN�1��w"[�e�TR砟/aZ���%_����Dy�!`:+B�w�J����^q��j(u��`��_�cף柊\�7��p|^�n��(u <��=
7��z��M,D�P�`1�x����ǣј���^x�����+�	@S��ؤ6M09^NĄ�<? ����Y"�k�������'XasҞ�ˁ����pzqL��b�9a�[CĐ��$:�m^�[c�fH>n���e<��a2` 3�׎,찭�U�v���."P��B�71�6zf�BgM����S����Cz���f��XxD�<��<{څ�ý��}�$��xJ���b��3ąX3Ţ��4
�55�CDH�Z����!��G�)F᧭���,#"G`*�H�Õ�7��#���b��Y���!P۳�Ό�/���a�/�pr&�4��?3G#�o�z��F{��6�fыIC;+~[a��{�of�U:��< �矠������C�qu�"�ZuZ.�Ǩb������I��?�����o`/�J�'qi�&��4�Ũ�%�|��S��q�Ķī�rN��{�F&�sQ�'��o4�Ā�N��x�8)�c�9��/t� 6�^�������4)�N�8��b�#��Dh7�t� -P0��z��8�Գ+�D�	��GִY/��|]lׂH_�^�@���0T:4��|0�S��D��?^�WђY�Y%\�F��xPj�L��΄iX���\��=|��!�ݜ�p%��#����Ey���<^��d�C����BG�0�פ���'r�C5�����I��軷
O+Z)�Rg�ΰ���zX��:V���ґ+��&�d2F�櫢�uo?$��r�(�"j� ��t����	_���1w�楼jU�=іD}e`qFn]Y7�f�I�?�
HB6e��zQ�t����_'�(�������F�!������;�d� x���3���,��N��2�r��k�{ه�K�1r�W���"���Q;t�2?��y!��LHU~�媃��CE��nn{��a��niv�R�-��O���Oz�6�� �!󼚬��|�8�}�,aJ�|�����~u��j�R$��L��z6� N������T�C��6�!y��ߵJ�mX_�8�u�&��%E��^�۝A�����"�v-/���;UT��N�toB	�JW2�̠J�Z�A8���Ų)������sIu�^�J���!i�Y��4(u�H%fN�~��!Sc��_���l�7�n�I@É��_n�����w��.^Ƨ�k���&���*%V�xp��c���h�aɟ�
jt�p'����%z~��,���TN�nrȴ��aGG�s0��Vz-��c��R����ܜ��<��Yp��o,��Ձ�^���Ir�z�&El�ed� �D@jgJ-��zJv>&\��t��1�\��	]��K�7���l��㳾�5��&���':�?8+ԋ���'��]c-�M �4��K�эb��h��3]�}o2�$�W1�5r/`8�%�3�w����ҟ�Iu��*���f`R�X~n쭏N��rm�&��&5��a�FW.������*�Q��B�.����Io�2��u�YoɖE��ta^�� J�"�G����9]��x�����p���z�M���"�/_^�����]ʈ�J��k��I
���b5S�ٌ�kck�I��X�yZ�s�+oY�O�h<������B}�ՠsHem�[�T��qS���tܴ�eUG%'�b�Y�
�HlSF��t��>l�8J�)�k��?@,�`hL�>�y=��ٽ���G�0����.�x%�.a��' )h��Rp�pLk���g�+P�X狤��*$���#ʗj_-t�Tq�?����?q�x�^*���NvľET�U���ŀ�Bĭ�0�h�GS�R�D�	�9���J%q�	�m�a!#�����ð~ �Qa+*���Н=���>�����@�١}_O��d��*R(�]�{;ҹ-yN��nX[��Jҍ�[ZAZa��B�0{ �א"�s޽�8�E�r�i��ث����?�&����`���b{����&&����!