XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s�C��v�l����h#��bjA�U_⩖�K��F�.+fo��D���-��я��Ȑ��?���<,����@]�JH/��D�6�A!��UJP��@���������N��X��
`>��k5]n�NK�������q�KU�6_s�E�%&�u��!a�?u~q�<4���H�bO�&�i���M(/8`�0]�#����m�\MzV�=��kO�K��y�apl�����-��W$8�y��aIV���b�#�Y�j�-I*��%��+����y�`�A����`�S��Mp��YO���4��1d^Ƶ�wCV�]��d��d����o�jC��׏?r4ԫlY!��7�����߾
��g2�t���a��*�,�1�(��S�0�s�  '�ii�"rݟL.V��l��&�!�Sy,�����j�`�UR$t���1W֒��EN����o<%��t����5#�Q����\�cOw:R�7�ȕ�N�R�G�W��=���2[��K�V��N��կ�X	XŽ�U�:�ۢ�8��̛;��t���>5�7�<�;*�l��Dd�g+�3���o��9ٌ������٥ 4|y��mȩA$+
�4�drX{��c�7p/��2�ߦSkcw��?��k=ȺYE��<�7���u�G�q2��R/�		P ���X���qq#����^#;`����`�M&M|Z;Qe�5�W}���h�Wa���t����~�g1k_��d�Z�ect�X�h��XlxVHYEB    fa00    1fd0����2 +�눏~���T3���m�2eP�Ʋ2��U�=�Ϲ���{2�Ѷ�#}ׅ�n1%��NCJ���`=Sv�t�r2�b����S�c�Ο��	�)��Y]��X\<�͑_������L��&
K�����TG�f�����D|��=콙n-���jđ�d/��� �5DW���.*�0�Yǃ��|М�n�k&%_BE+�(Hf��[�7%��M�co�x�KM
����_CP��%�*Xj��";�{���7;*�lSI-�v�*�~����oj4�S{-��Jk�ㅪ$]%��|�F@Opϫt��D��e|��RC5<����E[� ���#]W�YS>O1����'���1q��yCg�����Q�x�jV�X���ٰb>�7�]��[	�I���}�QE�VOm�֑�)���|�?N�Ţ�W)���2��^�K�X8��ک'��ӄDޓ$HZ�*����+�E���e��>ln��9�_J�	���L,��(qω#������;i�GC��f��q��v�v�7%rj���Y&'l�y\i���u}���Br��- ��/jls���I�o�P�&q&���p|1OF�bpW���a�)2E�]cbmY-!����>��m/bT1Ԣ����dp9����^щUnM*:������e�#/��6��=�9�V��"�r�]����;3�@�Kz��%B^�׎Q��KJ6a6��(�L�("�]��$�������[jO�<���S���U�|��:��#��ۑ�t~'���Ma�מ;@<x�X�������#�ب5��(B�$7�}��/k]�2T�#f��2l�Ԭ��܃r���p���-�Z%,�n>�"�X�����Y�o�L��"Տ�q�D�J�h���a��#`������(Y���q:xj�����&ɏuO3��H�U�P�����e0�Ҟ�S訧�;�)�d��L�.�)�"��?�]E!��UK��&o�T�r�j���b�G���Z!�Ꞛ�ǘ[�
��?³�;�\Բy��ʷ���h�zb�!���gk�֤�����c�h~ĭ>��V�T���WlU+c��๼l�k��^J�P�0�F\���6��d��T�gm���ׄ-�̱�O-/�ha�'f�U�aHr����ܵ�kb\
y"8A?�U�|v�Q�H�tUc1�,b�/�AQ͜A7B���q@��)�����K�q�h��|H������@i���,�>����$c�>T���K��j�x?>&�!O9ǳ�F���k��P� ���S��GF�5���� _O�q��Bn�/
�v9���Ch�����3�'���[h�S��!�A�d�I[�cC���4�A��g^�|���}��V6��5i*��{�qq�J.K�� �[��@��A��ƕ�4�G���:��Gi��h*��hD�K;ӣv{{���S&�F��kO�z���>�S�j�~�/���M�l17�w:Z���࿴�3���E��IJz$�PM�[`����S�������ߨ��B�!�|r�-d�k<b�&���u]��M�j�H5��8q��׋����]<"2�CB���A��PH��;��Gt��ׇ��K���I�v.����cyg���
I�����f�@b���/<a�Sj�Y�	���ا��^[������#Ldu�hK�x�XE7��g��N���������qUVO'E�������x��K�4���l|r����'�E�-��D�Ӝ~��m�^�`��U�SE�S�j�/�|�ق�2��۔)7�L���&�M��c�S3�y����������x�묌�#[%�>�o����۷�I�n.��]�A���dv����������~�*|���d��G���&3K�>Ħ���㕘ڙE	2T��/b#xub���9�J����T[��P���'c >�� [��	�Qi�	bF��֦w�"_$ S��(.�Ƥ�`d��D����R��vVXQ��/���9ub��K�4�k�Ҽ�F���;G9��чv߹�J�#2�2x��芳�]#a�5������a0 ��+��Z��<q˺o�=А0h��@&������x�P0�'է��V
��3^&`����2d��^S:'[F�2�
U[L�9�x��&2Q'�uPI�2��Φ�ｧ�%�3����KHC!� ��r�}�y`��j�$���%	����c�j'I�l���{���#��	��z�zJ�>]����A�g�a�	���>���Z���u�}���=�6�1�{��\�^Ήh��A���1~X������^�7�����qv@~&�e�[�]�C��2���"7���	�����<���2u�W8�	���6\�Eh{�
�]���pC�z2~�)H��<���t��6Bn�'a��E����-���.��S%֊ow��*���%�`.�DxH�����O�Y>�v3�J�-��d���,�.�z!LG���(~'Q�C6��fb�c1	���*~�ލ�?$j�H;\n�7Lr!�"Ϭ�������薏�Giֲ��hO��/�:�V˯C~/�Q���R���σ`�V7p��uFټ�&���Rwzn>�?�IT��e�W\LF�K��it`���p�>/�9I%�r�{��\��˗�df"ܕ�0��Mk>%��=�6v��ۄ��Qڎ��L���E#�y�Y�ҢfT�.5�dŮ$�>z�r��Dka�o�˰5�����h��U�Wuʎᩩ:��?�Ko�?{b�Ӌ�`���"_eu6>K}8ō�A�7���-@����߻x惞<'�����![�r9��kH�_�qUݩ�b�Y<*�'��ᖠ�J���_%W�r��Q�{�](�_!o�'�������Q�aC������5�� �s��ى.��Ϙ,Z1
?a�C���4�C/�=6Z���}@�4����I��9m��H�;n�����DE�}�i٭#Dqђ�w�pc/�HO�`���Z���Nr�r(�F�ܲ���ո�a�q��3^/��ln��Cn�����=��7�LZ���T�8%�ٱM&a��w��JxD���3����s���G;fn��Y��[��P���CPgG������.27O(q�A���J9�<@�t�/W���#�m��[Sּ�~DC/���hKv��vo��XY��z�r�qyWbrˀM�a�w�Sג��x��S�=�"j�7Л�����%��G����|���_�o�� ���R�<�]u,Q����1�3�+Sr�XRިY�St�I�>��W?A�t�8�w &�Ů��hF���$̮�eu��Q�2m�F�����>%}��!<^|���*�R~ڌ�L�G�����Ζq�F���$�U�y����S8��(��#>����b�^4�}� �9ۘ�]��fh11��5Z������/�c�}TЇ?����q�mPV.O�E�G�����Ix�;A��1�|�r�a�����#��V�*��'�qH,y�?�IlOl���F=�/h����5J���L R&k,���D@�/ǋ8�z�͏��G}��Q��y���?�[�Z�WO�<����6�U[f�=@�Bs�>0�5�����#��3���b���d��D�Q�H�4^;��8��M�`���s�_fGW��	��J�a���Qg��$�v�S���_	�`�=�������EY*[���/����t���BP�>l�r���)�
�f���*�l�H e!-�IF̓sy��Oe�V=�D,�>�����ڼ�e6�i���N�{C3}�-T���pxC��������1�����%����o�|K70=���L�-��-���!���aR����<W<h�m�q���~S��)���=�}�0�l�IR��Tc��AD���2_�t�y	�cp�����Ǳ,���PZ:ui�P��5��#���8�j��J��[P_���ǸKj2�g���,h$�f4�-4qC��xQo��OG����[��T�h�	�����t[K�/Y�b�-vihE�F�����vWI0C�_�0����AJ����8^څɺ�mI3��R#�D.@*ytug��R\Z{ڣ�ђTx��r����U�gdʙ�p�sh��:""V�6&}����%+��`΁J�g�Q�tKߺ̥�'�q;ۘX =>\�I���F"y4v\6�/�4���|���lU�L�i=G��f �&��@cÀb,���3��������cw0�D.�����zD����ú�B�i��o��dR��BD��<���~TP����D>a�[�G0��(Ś���z����,�I���픘�B�B]�N_z�8dKr b5^���U�B�w��g~������w�F���P/j�.i:w�7�D�J�S��kH�}�8{��>� t��B�)��jтo;YW��#�I��'�~�֬8��"3a��c�1��Œ�d�e��B�	���U����
~��	��Q�!a��>������_4�>	SQ��E �==8�i�B����j�WU觭Ɂ�-Q�z�,���)���:�U��yt�ïc(�.7��]�6Ee�����y/���ة��C&��Ϡ-C^����<Z��|mhZӡ�BJ�<�H=�"yU�~� ������w��Z���DJ57~���Q�./�G��2z�)�w+�(L����r&�	���fn�����s��t��o���S'�:X��^��ŗ�V�{�lw���y�U�>�Z�?����_�tÙ���/��W��	���KT�3g�Y���iH��X� �t$�x�̮�b��~_ή�ؗ�bH��^�
A-5JV���vEa�B�,�uD�qb�`��n��<���7�˒�uQa�G���X�gԶr�����~A�X@����
UkT�L$���2�Oi!Ӟ<���~��_K�jr+�p����ګ�_����;����9+l����H8�C�\�P�cK�]�e$u�r-y�)��.#"�+�җ_"g��lA[�O?-�Tҷ=1�Q���l�L�2X�a�p�e�-9�L�%:.(�J��$�4��5��\}9IQ�/~�у��4Ϯ�E��_t�+}4)��y�4�Y�@F��W�-�}�<�R�L�||�܆x�@�
�7���/lk+Z�M�PA�;���0�LL\)��R��}�ch�	��RW�JI�B1����V���e$	2R�6�R���έ*W��}u�vP���H���){wC��^��d�����}�b%����?��	��:�R�#	{o߇@�q��u~<�@3F3�lŏU�ʩ�y��)��-���0�yj��J��՝���$W]3sYH�Ͼ�Ӽ��pa�$ /b%�������Q����΂���/�,R�ͮ�V�<�h0�e����#�l9��V��9@�f���b��UI���q���y�%!'e�1?2w�D�[�i\��(���մ��ɿؕ��n͐/�ˠ��K��S#VwḚ��)�)��5ҭ��Uv�'l�LK �������c�.�ks;Q��z�ķ/{�4��º:]��wkx°aKD�5B�2��x2ƁPX���Z��1�	hW���?����,q
�����B�j!1�m�t�s},���,'/Q��L��>�I=ѥ���K�?���`�nF����+FWq������W~�ku�����7u8b�(���8�{UH'��p�"ú�]�j����+4OL�����p���Y��vq�Y�K��@W�0���<�1���dZ������B,2BAY��̶���;X;��VӊL�y�����踇NH�_�=۪��I�b��������[&���/�pdъ qDP�{��NH!�i=��I��*���n �	����UĕC@�*�L��#�B������*P�-����;�M]��I�-{��6�p����Ok�UQ<[O3IKlz��� �$P�?~��l�
�*õ"�l�`�L����՝����e?C�w����hãh�9����XnN����X�i��2d05W��}�!�	S�][�@�9�y"m8�E���nڡ��Ʒ$Z��q=�F5��n��bUҥX&��d�i�+�I�.�d=����<)%OUnO�/���/�n9��~��O��J�Ӝ�	�[��z�"B=������;Ky�Y�Ou8m�$g,d�&q�n[a5�K%���u���˺�͜�l6ּ�j�Q�4jt���X��a��%I�U2���Ogd���bW�r7���p�{��"�r�-*I���=7��$��Y���C�T�Hw��W�o�lb��P���;�LUJ�9��ZG
u:^(n�S{^�u��[�	J�}Mѯ�?�g}�?u����K�)����os	J|��g�f�^ P�{\D@c���W�j�9T�&&���~k�+i�>Nr������3���ss>GU`.�oF� J�3�&v(R;�1�ֆ����}�����:�j��͎X�9k"��Y�����&�7�W�J�$n�%���lWsC�-��=��Y�4�:����/uJh���L:��o�x֐�@��ѧ� $w�nVm�2�yp/Ǻ�`��F��.�s�n ��χ���]2�#���2�d �t<WA�ꒈĕ;g8sVm�cv��T�J7��o�= ��U�.,^F�z��]��ɥ9:F)XD�6�KdK�]o?DJN.�֡R�a��p�b��P�����-M!��M��c�k5`G����#5�n����ۋ:�N�E����Ȯ!@ !���s��ı�I�T�v�4�%��Cq����-��ͶU����:�� Y1o��0�Ci��"�T�����Tm_�l�:ǽ��D����݅�!�G��ix:��c��������"�\N e$��[�@��v1,H�yk�+m&��$�Y�c��k�&O�L$�K.����KI�Ό�oS�(��z�M�m;;�{,�Wέ�$-ĩ*���,7?){^k��I�{�J!�%G��O�K~_,�L5�4�2ԦU�[��N���X��������0�#%���Ul �8Zj@����d��/	ᴤ~�ә�V��g-�H�>�/y�����:�|i'���Ί��� *<��u���U#�r����z���)t �AЯj��Cs�oj����ܙ�
 a�^��$�.�{`HzQ�}��S/$W'��� ��-�����st�ʶ����)��2ʪu�^0h�h�"r��0��"�(}kCt����ob?���.���i��ՐU4p�($FКr�E¿�v���LUX�ho��W֥U� ]���Rp����oP���g�N�L����C�������Q_���!�+a�/���>f�?Mq'pQ)�:]m���(��4�Ϙ���*8�¹�_�W�B�[X6@��^��}���><�2l�&�yc�19�xݡC#�8!��)Y����cPLt�����ƌaR j0)MT'�� ���~�����Sě6�#	�}�g�L����"
e�ٌM��A��h��[�!&�,��w���"��;��K�n�Ǝ��Ot�g������&_��K	�X1�0���
$�a�m^&�<+F���T�<�sS������Թ�C�H�O��Ͳ��QC��f_�B��PV��^2(����!bU>��jP�c�Z�� �! ���Z�]��šV ���~H;�X�A|Y�AiL�כ8��<�X����p�Ӵ1"!��������'%�z�S���ƫkf=�8�|DYӯ��vsW��~L���[s��j��={�V�QS��g����Cԧ�Z7���)�?9(t�:&d�S�K�|]J�L�a��h�lNWF]���(Q�ʋ֖������&���s?���`πE"����)ȿ6��TpCn~�"ႍ�~U� a��)���ߵ�+�h0�\�jb��J(�@��JWh)�P �Jg�[	��ŉ�Y�FGB��A�a�n���ͩ�(,A��]T�V��C��P@Hb����)�\��\���@|��vW
�#1?�s���Uh�R�=�a�&#�����"�XlxVHYEB    fa00    1340'�4U�BP���<4k��� ��������-J���mS?�������r�z)�嘦7�T��i�9ڦ1���>z|u.2M�tD��3�&��6�f���ybjT[Ѡ����h����5>ҧ�x6��eiq����	�z�IV����t�I�B���6����e��<�g�ȰK���wo��G�� �Y]S�2�;T(wH��-P(�{��`2�/[!��3G�t�!��r���@r���2���Ὠ~�W��"wFB.[v�̛����`Jp#��>$��`��j�����Ǟ����;�y$ˌ�k'6!�k��(�˶C����l0����uk�d���G�f���[6���p���K��<���>|Ҵ�0L�Q��uC���<�@�$Vp�#}"3���Ѭk��0�?����d��F:�,,(l�!��ׯ�/?؋�c�܇)渹+ɅWV���͍GX'u�R�����vu�{>�N�ɩ����\m�!#����-��tfHD���#�I��`�NFp�
��V�4���;^r�hy9�R��dm�T�[�z£@��쿦����?>t��s*���;]fG8�X���|`=?��]�nي�:�M�Cc��gJ��`�:Źb����?�������^�W��b�DA�4і,����94�(!��,F���:�$tl0���Q<��2d9Y˗��a�M!!4�٨:�-c���Q��t�!�6a��k1OΐV�[��MGj�S\Be�&Ai��.$�]�"xO��#������p"�|�.p"��e"����qX4��ٞ"���"��Ӽ���a�>\���/>)��J�Ir����xr���/C�tDo�I�Z��UB9��2�	�8��fף�zYJ��VjM�O���|�N������Y<*\?���*�~�ũ�����ܭ��!e�aGT;Ej�QE�Z=������7�W.tG"2� X!$�T�^��ۂ�ǳ�R�`�IN;��#*�ev�0OH�gZv 
���ͅOڒ`�5Hv'��o>���(� �
��$��b?����e6�1ф4��da�Y��Dd�����9��:��9��6�O�A&{\�a]� l/��MD��*8�zEȚ�l�"��;_�]�A!��}?���Vl�-��dny~˩"(�q�$4X���0�Yl�9)!"������N�C��y}�m㮉k���
0k���j��<�b�������b�E�v��W�/��;)B샜�*uX�<�)�vh����p�Cr�"��Ca
�x�x������xsK{�S�BI�w��ܼ+�j"��V��kl�uJ=���YErǯ_�g�Y�1g�^��#�5C4] �>��y���߁Jȼ��W}��B���B1S�����8�xĢ�@l���w��e����x��W)X���2�q��%$k��X�L���)�M:�>a� �E���;��VS�2ި�G
����'ٙS�;��.бu7'ȿ���q��<��I��豆��y�q��;���.0�
�9v��1��Iha<�7Me��ܥ��z�c��j�A����������9� !L�g�đ�kUD.���^�j@s��%`e�y�B��ɚ����|�lM�� �Oi6/�I��d1'�ũ�����AA��+"��#+D\s�7�rtv�^�mr��Z>�h&�*�!*R��c�EM�܁aQ˳9���߰͝�����dE��
�r��Mx:G[���,�l6��C�YkCxA_�}�#'�c{6���@6�b�O=�~�O���L)B�@�$q�Փp	)&O? �����^K���!3#��"W�}����m�]���M��WOJ,��pf�v��!;)V	����"u�?	�>C!ZT�'kF-7�}���g�hLig�kmj�i�A�6�f����O 3	vǄ��������.���1������SQ&��L�KJ�$��$)���c 8��ƅϚ� _}Q$T�/�XC&��7���������*��E��g�����q�[j�߇�U0PQ-�@q^��#�Hj�˜���sr���V�iU���ӓ�6 zrȣ��
%S�P�_�A:��)d35�̇tO���l)�#���ֶ���X�=��LG��E,C��g��K�Z��oZ�Bo��@K�d���4v��R���$l�����O{v���:Dg\�c0��kǁXC!��+�;�Pr�5Ԝ�P�@����J���|��Qdp��swִw�����m�{�f�g��ԏƛR=�Lz�
�(�������!2d&;���>xs�g�t�9��F�n�348�FB,P/R(�a��}����+��֖D o���JL�)���p�W�T�E�AYHͣ���ٳ6��\_�I���bv��3x��5&��侇���}1�SR�Q\��׆����ݪ'�1.Zrh���Gn �Db�n�/F�|�Y$߄�E]�SӦ'$�i�Q��g,�����i%�y�lKȏ"fM��u����DKUb}S]�#�Ƭ��r]w�o��͹櫻8-t��2��_QS���R��qr��`#���64C�0�Ckۚ�0�,�jp��Ro�G�zI�8i��%�F�b3	��y���9}�\�i�g��p�8OdY�#�_ԧvz0 WR6Cf��Y�Pҽ;�����婠&bH������;}� \>6P����sX~���)�;#	ũpk�ԫ��j�S�؃�/�f�'��m�7[?Knkf��g�ff��tΎ[s���P��^�տL��2F�����蚍��N'F�J���brYT���6Un�l{c៤�.�HB��S!Ab��)焕��!�����l�:V�i��&Ά��f������F
l$�-Ѽ��ނ\�>���]�׊�]�l��<�h N�s '[��x� һ4l���H��{��Ѝ1u�dy�/D���|���ZTF/{y
ݯ��xPě)8+����5U,o����(b?l�m�T�!hb�Ѓ�=�˗��t 0O �nIn�n	��ɶ59�?t�bB�stP��My]M���]�&�%[75}n�Pd`�iN����1;��T��`�$4w�C��@wx�_s3��d�qa�S�^�RQ,W�s� �xAk�6�I��s��`F����=���}	���W�uk�6﷬�5wm/�f@���kC~����<yOIe���eS�ſ<���:���ؿ7��`.���y.FR�{���u��1p�K�'<���A��3�Q������o9P�-k'����~�����G�=�t��
����i��8P�N\˲+E)ɏ��G�㭃\�禹ҠaK�(�Y�s�&|#��x)�rt�E�m-?!�Kkfl�ݲJ����ފ��O�wg0���qi����W��K"��J{�=��٘�|���[2��ݒY��#���%Z�,������G�}�W�M��!������H@��%� �MsnW�OkBp�Hy��.��DdR��cU)��Z�gl�MM���%U�A�E�]ˬך<�w�`]�*rQyN�m���j���$�枽Q��#(_z��l"0jJ����%��6�o�_��x{D�3��t��۴������/n�c���CBOmnZ�Q��Ҹ�o��rr�%x��ޣR�)�$>�bI��-�:;?�N9\����7|'ĬnZ�{�ѡ!����_��_a�'&��1�?g����h�5���'�bf�A�x��paBl�=M+w֮J�t m���Pq�� ���d)�^��o2\b���b�@��_��K����8���t�{�,^fJvy�V��?��02���T`������=B�5��{�}ْ�P��󕺰�B`#�����j��ԭ/�[�<<�z�q�V�-�Xu�b��Y���)�bMc�G!�����2��h�̥Z�T�G��u�1�F�sB�2!�j�J!�2E���v�K>$Jìڨh�L�h�F�oiq��������N�[���Fڼ��Kq��L��R}��BB�q4��</n��5�	O؈^��+�fjJ6�D�mBMjľ�p��TKmMk����5�;���m�N�.|�c{��	�F�`���ե5���=���Y;MĨ��T�ﱭ��yY��<��-k�H�0|��2���7s�"v�u��N�+���Tw:�n�S
��$�����1��y�:�z��4A�ٗ�5�e�m��s����3;���F{����k~�
L��TU�i��@|�wy�&=�.td�䋻���#ޣ����� C 1}�� ��~T�K�P�n��(^��Dx��V$������K�0J��\���I.뀟�ܮwm3�����2	v�M�^"pyT��C�v�3��C`��w��	�4R�l���y?�5��� �9�e:@����鈛�T/�u���ʵBx,w�>yG�ؕ���k�	&�~M���:J��"�3��j�-�Nꚋo5�S����'`����V�F�����i{<x1��'�Tf�s��C�����Ù��%S�\�ao|/�>5,u=_��\��;,�� b�?����2!��.�r1�Y%a����9�,�~lT&�,�s�tH��P���OZ�?pXZ��������my��PP�~���ӈ����D�9@A}�����e�^�U����]h���6�Y�#�\�j|�EF�����i�Vj�JCe%*�l��K�C�P1�ɪ(f.�h�]|9��;�r���A��Ơ"j�k��K!��B,�Vb/���H3�~�(îHB��U��{	B�'d��
c���q��^�Vz�!���������~N�u�\��/`9q`+�,���s]�������0���z�K�?��XlxVHYEB      e7      a0��`pW| ���<�:�q�����ڹ+�/D�Ԫ�5�koJO����p�Q�{�?q��f�#^$M����;��-*^#Τ���i��I�R:((�����Z51韮b��i3����#�Տ*~Kjrc+\Y�u�Л9�N,{����zb���x!