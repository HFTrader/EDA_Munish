XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����5��?�X��
�:�B�zd5eK.[��a��;��N$]�����$�D��2p	_#���?�u�֣]�v�kR"�Y%�����+*�����iel���-�~�>�@�����W�h�+*Lu�x��JÐF``�{[�:d	@���c�(�Al�}�K�J
��*%�I�PZz��nzͣ�� (- :8��֦������#,Cg�^�5L�պ�A��M�i��\��E�u���QeY��WXЙW����4U�/=�sF5[�w�k
 �~�a�@q��Ng�8[:��w�Q��t��[q���zp�H�H��2:�1�T>�W�*��H<�F�)<���������:�٪��u�3ʻ�o�cun����
S��Ǥ�3X��c�iG"j��Q{UQxmQڱni���p�aK@V�R��0�3�b�%>����I$7|�9�Ǧb�IW)��;)�9��!��y%�	��:\��q�����!#������	�����&�Is��d��0��Ԝ7VcsV��~XĤ�A�Oʬ�*�$"Z�B��m�q��~f��� �m�r��h��᪽�Z�݊�J�֣�c�׍g��`�1���G��'�����qlH��X�1X^��D;� ̇�~���=�ߦڳ��o0��L��ƾ]�����Q=u���Yʢ�����a�z��l6�.X��^u&���bgHNOНB�R�{WIۣ��'��vf���������DU`=f�0��PXlxVHYEB    302e     c70����e��suȄJ	��?��� ���O^-I$w�w���'q~g!z�ޭ`��pC:b�ziϓoT� y�R�PK��a��Za!�G
�MX���.(��I�E=���f�O2�݅��h�!t�pj�)x�-k(��J�8��p�7�s'��7\M	���,��ZB)l�شk���	�&�8�kia�Q?�X׈�@;����@t���M��H/���p�E�#����2a��+��� ��r�}'sjt�=�Yܚ=`������XV�72$kK-��cS�����鉸�%=�N�����]tU�ʫ�W�5s�[��$2��_0:��c~pO�1t
�̃Jہ�&���O<R�EK��1d=�ZB�!z��VQ[`9dre<u���{�ᵕ%L��a��9;��j�ac��)���h���[9�*(%�!Fi����	+8�)�4��S�Ҋ��-h��~P_���۳iKq�dW����!5);���~k��!�e�2�c�K�vI��޳i���Ҝ��2�B��PL�'I�����$}�<xo�h�P�z>r�w����(��z��p�;���Z��'�k}�f��O� J�X
Љ�QO�J6`���zӫn�^-�h�a6�az&�,�h����8CM-�-��nm�˰ TE�����!��2�3��mw�P������0WBٍm���-�J��e�!1��3qC� ���݌v9T�l���r��ڰh(��L׃�WC��;i�-f���o��M�j��P���17�~�%=�Ȥs���v�P�4MSv:�z��BoX{,��w0�����T���k\#4�\����-���!Њ{��i}���#CD��yMz}�I�W�z��P�G�%%:�L�ĺ�@NE`$��R��Ɵȴd�ӝ��`���팈�;�k�>�,f|����bG��:��ʻ����$�lu{��[j�sf]���1�zc�q�{�4�u�dҸwC��<�if���A�xB��Y7��B��<y$)-.k1�7!t���!1�M�Z��8��=��q����4��ou��M�*NA���ţ)��|q�dԀD��\��aU��֒����)�`����2�J�����%+)ߚ���U����7��t��F����c��`���l[�7�K� �����*çp��L#��=�7+�Ox@�ƣ�ŁQ�}�[yO�@�#���)���.V���Bw���j�@g�e�U��$��sƒH���W�)_�m]!���$_�����ȥ��x�����zT*	u�7O����9��H�įv�������g<R�徑2���y0�#�S�\�wy��ID����9���F��퐴�aįDľ���3* ��L�,:���4�"H���I�	���j����wdi���2�|�Vt륚���b~zQyR��a�%3A�=�jH��B[m<r^`=�e�E�1�~�\D���Ӧ�}�j@�J��}f>X}��b L�1u���m���)֜�r\�&1�գ�U���]�-qv8������:�O�M��ȡ�A?��E`����<Kemł�����m�J�F���4q�;��x�	b;X��Xdk�L�/+�E�IG�j�]m��z�K��i�[�U��&#v< ��T4ӢwN��C��R��iGL���)K�������P}Z�/���zP�-h�4dq_]���݇�HU�J��Xs��.;����ƪ��n�->K������^��T]&^ӬH�ImA��)y�!XQpĎf�2�c�a���A����^$9���������>f��;=p_���ý�
<j_�S�s>�<\��W�״-j�I��CEGmr'��ه�\�K�~��� 	��ȱ|�A��fҶ�_������7�[��'���w���N�NK�k3�'0ÒG�fPp� ��{��_7]���k�$+-�� �~m��_�}��! �[RQ~���j�j4�4h<CT���"6G�����X^�q�����W����t#:t]�;�)VU��BA�4>����L2t��� |��/�UT�kT�K,Ԓ��P�����bǐ?�Y�9Jm.�˃��`| &��f�P� � ���!���(=����m�pZ��ɱ�r?�'���Ύ��(y�C.����ѩR�8}����+��VzQ��r���<5x��@<t(\jr�ǝ]�Uz��Ęl~�8��>n��,f�\$��@x.�N��P}����(]'�[!�/GU��:����ݷ\b?1@�U��(�;��y��x���y��}�fO��e�;�����^����j�X�4E�ٴXs���VK4�y�ہ��Ed���J�
�!M��a��m��4�y1eo���c�[�K�?K0��x����m�`
�Ú̮�]u���1�ڣ���чj��*�hu�Ed.;E�}�� l8��~�:��'�ŭU	��B��|`�ys��7�����Ϸ��1S�$m؋=���]�n�u!s��m�ή{���6-@���>p�* �|��υ�)�u�,�[��K�a����\
~-��4�G�}ع�Z���Ar#�6|����j� ��.�9�"�iV��f<@� 1I��h�T�u������z:D�~���a����o�K���L��t5�oA{��H?K�ހk��tEZ[mb��6��.�Ȉ�Ax'�k)��R@R-�/����0��Uc�A�5��?�y�@�`����m#%a��+z[��h���R���Ro�T7t�$$re{X�G��+�	|M�9���cs�2&�m�i��;gMA���ZOCχ��x#w���%�T��P%�W���.a����0'���*����>p�!!��Nxџ� ��I�a,X�`��O����6��qz,��7��N@�� �e	b~��kz���IZt�ܡ�B@�U@җh��$��>]o#"%m�������Sj�7A-G�.�q�z�+}x�UHL�+�y��s*��y5wٺ�v���딡#�r�k�tC�����oP2������2�%��������kG�zD��k]v>rBBok��<*\g宥�a�_X��c��@vצ˄���э��*h�|Z��de�h�e���EU�%T��B���#���E�_a{���>%���S5K_�3.sW�?3q�w_�m���9