XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�&�|Z�PITд��[��O�}R����Kᅴ� 1S�=���X_������c�Q���s�oX����"N�����ެ��� F@0�>�hn�{�my}ρI',="���)��b0Ir�R��y�a'x���^��6II8[&E�RX��Q�A���I7RQ&r� �h�f�#�o�A}^_J��NDCd��ИDAS��tV�=O�Z�Gao�_�{�0wu�r�"�~N�r��1����p�9��dR94�:����l�D����~�f�-�	�.��-���w������p	�\�b
� ���$�ku�M���%<X�������e�6(�bӯeʤY2u���\5����l���P�qTN��b^9NSΞ�UK�����_�ZxY4\�yi�zO���!�;䡬T}��X~w�1i��՘�}�����tlI�w�����+`g�g��=���r���R����"ҰiX�-2q�LIaBM
�}��Xpp� T`���U� }Qϻ��rn�iCS��8O����2(U����h0�F��������si��=*3	1��%����J��P[����F����ۄ�j�}H��bv���f�u�^rFK��t�G^�X8M]�Xe�]]k�k���*�46��[y��e��)8�d�jj�.�*{_^�!6��,�x�Q���R�HI"�=p��9�#k	BbO�F�P�(��Du1�(TI_���l�^7���K_9X�Z)�ܽ�HR�<��"�XlxVHYEB    2533     b00^�<ӏ
��ת��������0#v��uP	��o/vG%��o7���V��"��k~ ��ۏK�~���4l)�$*�_gt�f����>o�.�l��W��B���Y'w�M1qK�YJ9��h~��X�J���rTa.���W&���e2�Ÿ�s3��v/��8��@�S:+���ء[��S����
?�6`mg �[Z�/�ǑO�wS۲Pʿ���1�(T��U`��4���N-�#,]�y�q= ����i!8)��f6r���bm:�>�z$�l��f��֌4L����%Cw�{WY�Pb��]X�j��k�c���L�$�t �5)�+|�Fq'�>�5a�#���%yՙ��IJg~�"G��X�~ǻ��p-Rcm-�����4��Pm�ţƓ$�\�pk2S+ԍF������
���.�>���>�g���S���Wi��ֵ��#D�hY0:B��N��e�����M�j]��a�(5c�-�V{|�D&��^����|��!č��H��$���>����D{��(���=�.�/X�O��Y��岓���b]F7+L��Z����������Up(�g�m����(c6�NBOڕ8�
�&�ā߾҂S�~�+LBk��E?	 R+򚣀\��C�) ����>O�F�q����~!hmWHZ���]x9�R(Ҩ��
�7��4n�S(	�cN��n��NtϝZ��Ȓ�ť%���?-ώ�Da�����c"�=y���Dt���H�(B����_�4h�np����n<=������#���dgX�3��S��o��Y�� ��V�����^���QK*�R��Js�X��a.A1��o>���t@*?~�6�����?�q����A1�}�1��:���ȍ<@A�p���*!�Ҁ���5��Z��*�
�$K�{�L�ͷ����OP��tRNph�$����*鸉k�.��M�-{n��>N4�X#��[v�&N����"�a4�q�m��?���h�F���j��*}5��G���D ��Lt����`�(*�i��u� ����A	�q���О2��w_��Etn3� l	%e�M�K�yگ���%���34�iV�\�� c˩�z�a_�Փ���hB���o�<.'h�"�exd���M��[=��5�|�tO2�SNiG%+wr/�+)�6��֮V��)78.�؝%�@M�H+ C�V���5�7~F��"��X���"�b�s^苺��4�p&M�K�_���|ΖUs:�X|[�A�8Ѳ����RL����SL�)�f���{ܡ]�u�x�̎�0Ύ��hM9�����hD�ڨ����q�8K~<�+&�7Q(���Pt^��|?�G�tmT��R���]�H��j��d�2�/�?�k�K�[�A{������i{/yP�h��F�^!	�jp	'�N��#[�G ��ԇ9.��n��>!��U-ZJG(�bỲ�wUe.ة�Wjv�ɱ��%	D��L��&}:��<��xb%�Y�î�U���4Fϖv���$��aP�1S�����vc��0%�����Z�=��Գ���q�S��m�ə����s��ՙooD���ذ�U��� �guv�p&����yNp���l��6mm�׹��D\��ܐ��+�Kȯ/���݄�&L	��Ji�$��ܤI�݀����d�JŇ�Et��:�h��7��,#!&�ˠ��l�d���>P�f\�����c+�2���ۿ���+kb$�5���sI
P<�:Ց��Q��V׹��<ec{�[%I�	�X����I���d�HH\�~�]f=�_]�^Rj�\gE��?bM��#��ؕj.����C
@�Owf;/�i���"S'/+%�#�"ގ���IX�&W�=�N��PK�f
aR�'��1|ļ�;�>G:�F�@vSG����1&��*[9|ͤ�N���9gV�]��{��Q�l7*��$y�Y-sEH�W܊dBP�
b7ݽ��T�4���Gj®�A[�^���f��I�̑��4X�[���@���j��/@U�!M���3�gcm��(P��g�`���[��:���NAai0֔��"����͜&w �w5�Q�V��` ����CeMfY0;!y�4�ҵ�3��M�^�B�4���c�,_b�o�X]�4��?�X�z�Aoo�1 2��ų���2�v
p{;/B�����9<��3��P�C�׵c���a�Zp��"MTؾ�!W���i���I�'s׋8K���%xj�	�W��ơ1)&��0��g=�SN�.���1��X����Om_� ���,�?bQ8�C)Ձ4h��r�l��;a��P#��^�0�U��z�y���j���l}��F��I����x�~cT	�%��.3y������Y��![�P����������Տf��:0x�/��6�X�Z#:��+RܹV:�Y �GCYsf�P��A�+B������U��h��m ~?U($�r9�Ep6 v���42z�jqz`�U�ty*d˄��'_���A�Y������Ye�P���f����q
��NGWj?5����-�|P rA�� �����u�B �͝��9�|"A2��mD*�-�R�o	��G��!�f	�
�$�Q��g�_��A�_��cFshO�x�<��ъo�t6jo�^�B+�j��T�����z���4�j� �m��\ǜ��}V�S�!�ܻ�}�J*.n��'Q%#��sj_�-挪B !i~���E�Ӻ��C�zj U'Sk