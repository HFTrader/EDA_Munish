XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��*[� T�W���L���M���w��P�����)�ô��y�$gz	c\��t�Ԛ�E�<,��@�'����Tc�?,F@�UJH��C[��+�}[�Q˫��C֗����2����ոV���=�A~1�
C{��`����ٴ�S����:8>��sd�,F�h;K�s^<r�X���O4�r��6��ܕ��J����Ѣ��T��¶��g(��L���>��4���荔�h����tSJ}G�
u�����0x���s�)�W�6R��D��ѓiݭ�}ǰ� ��{J�߱ӂu�����${ C�m=�}��j��0HQ�����f]�#}^����S�_̻%0��]0�e�1�`@�б͵��`	�\�<�D�Ԑ1��iV�4����
�O�N?ey�pt,���b�~G�$[�F�)?&�p, le}hO�"���N:ȣ�{�+�l�lsO�S��"������}qz��$K�?Q5@�/e�T���=��:ݫ�/��"I/2��ɖ�{
��$�/��>O4���e��І� �Ǽ�.�A�zU2���ї[8��͛y�
�M5q�� �`���a'M~�r�5����j��q-��9�߫-��g/��b�RY/�wc��p������[���ﮒb0RX�WiV�陃����w��,Z{��k�e�\���8.�2�d�?2�뛜��ӎ?���g�d��������������9+!lbt�������_�/�V�i�S��XlxVHYEB    2e20     b40��̓W�2(�7��{�FM��aƳM7e�&\�)���]Y�����<��1,ʡ�2�Z������O�
p
H-�Ԙ`8{�sOhF�e�
�Ƀß��<u���/�V�Y���;r�-�o6���M_2:������d���(���]��j��,�ީ��k��뷛
}�8�Au|�@�w>v�>��:WG 8�'���Ծׂʍ����O�ɲ�}U%R���k��ddH�3���ecѭ�Y�C�JE�/��xq@�h}Zq1�2�U:@*$ӈG���É�<��E넴H=�
��bG���JS�)ǏȚ�{�ct�j�q�`�A֍��E��k��'�k�|N�m�"� �n�nK�Y�Zr&���]1���N&�w?�a��)��ME����5%&�Y*Ӫ8H
� ���}-����>�[�|ji<�گ��gXQ��F�ϡ���`��b}ط.�ǃ�hDM`M��P#�G;���/եK����^�$w~12�	��A"��~�Q��U��m�c���{NS���p��Lr��j�K�Kk.{�"����H���� Z�D4b	F���R�?#�^�is�LJ�*s��b���e�#F���#4B���5nl����� �����6t͸�ɲ�I�4��6G sړ��>���p0t�?JW-��w�,_L#��j���r=�m�a8,d�Z
�7��hi��nru`�T?��"a�$��ޔ��� ��\��>Ŗef(0!;��O��c���Z���Z��س#�c.z�8$S�g�H��Z�^aj���'����@Ⱥ�h"lS�'�̳����w�pi��7\J���'�@��iv����I~�gT���w
�ɋ��e���t�&0��"�E.}�(�[�(�:��� �(<�2�R�ĻWD{V�	w�v�?B&tiݚV�\��79�ǢԷb�Y��u�FJa��&�K�$�9����:�9+�e	b�t-Xк�s7��g!�]$?���О��ӄ������3q3�� ćڹ�ڦL#���G;�H:O�%��p���~c�uӲ�ۍ��S�i�z�'��<~>'z/��^�mNvC��%����>��Yp ez�W�q8p�AT���,7;l�7�^�C^�� 1)�981{)O+�w�>�����1g�%�WKvr줤&����	���\�g�������§q�^s��9�j��l���U��?!w��aH�L�;��`�7�F�9l8m��N�
ݞ@T7�f�����\��7A�EK�O�T�!&���͹��Ly_8�㍢����� ��-���ѯ�"Y<h*'vTh2ݞ��
���vXD�;B�s�VDm���mPX��}�e�ҔDN?Q|�8�IjZWj���C(< m���z��p.�)�����������6����$�\�	%��\Qg���	ԃ,g!WVjx��'��z��|���F:ޞ�/�'7�qA���s�Pz�"�������W)U�WQ"Ɏ5>��8�\�hA˿Y
<��?5���H��Lz�	^1�����?���wP|7cܪ��Q�2��ʫ��5�/�m�˧�i޷�ﻷ��\&QS���U̺�����1� u���9�*��;gp�Z=�W^�:�jG�p��St5j�6�T����ʡ̈O¯���%~h
���ߔ7(�21�ǣb� y ����������Aϵ�p�����6q.ξ�Q�D��;o����*i$Xv38�C-�m!�/�~'W�7�]f�M�U]�+�]S���� ���D3Q�׼�Ģ���W�#1&3a�c%[S��i� �_q�ق��~KQ��Z�T���^�������؇���c�ԡ}��$����Z��
p%�BPD��gB��Г�ЮE�H�B��N��!׶^���nv��Tm���A�1�S�c3��M���P�#��x2j�2[!����Z�Pv��}0�كw���#\Sz�tcy���\��`]�[U�!�)�Dr5�c�8��b>����t��_n��N�Q������e���M�S��T�>`P����R�����y*0�V�� Bԙ��n�
�������_I�fz���}���(�}]��(7fX9� �;n5�������?	�A��k��c(��J��x� ++���\TzK�o0G��g�o�¥���0[yt��0�۸T�z�A}L0>JJ@��X2������H=����݆T!2N�lG����&�g igr>�^���Gi�ނ41)��,�"Q�cWU��\|e�x|�u�~ �VE����7*u�jF�j�t�ē�i��7"<�^z���S�&�d#��SMs�ߺ$�m}�%/�=���\��P��S�`coֶNQM�2����l��ܕG`�[#���Xf��dN�o0����4`(*�����5A�Щ<Q��P�q'��fo���()h
fQ�>Z����V>��E���C�V"�)֨Cwb��#��g�j��<r���]����#;R�h+�b1p
Q,[(6�S�ٻ�Q��i�T�22�3�]�v�2���v�(��E��	��N]�v�Pmv�&�I&W�o׬��z��B2@��$tE�_�.RB�C��F,�ȼ�r'������"���/��3.��;Es�@s��/h��K'+���j���y.�e�eS&�*�3����m���9�ݝ�6�"�An�6R�'oԞ��ul���3�v���{|�.��dqm��p�';�߅/�Ĉ�7�{Us��HpJ(zzX�.�c@*��Ę�Fu	��%� �gs���L���@�L��Y��i��z�r#���B��_VJZ�/�Dk�F�����c"����l-�(�D[���K