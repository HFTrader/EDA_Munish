XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����n"��GVa���"5~�3�o��*����Lc��+aAמ묓�	��������:u6`$FB��g�r?���NAֻ{~�������]�v��+#�t���b9���NEF��}5�q\�ڤ knj�0�0x��T�� �p%>ؿ/x�K��6�2��=�t���X��_|�۩CJ�y r*�(���J��z��3��c4:���H�q���*����#�Ĩ�e�|��:�U,���q+ʌ���BH����vE��Sd��W�����b5V=Fs�{������TꟗT}Q]�Yq�%G��@60�����M-�3�1'���` 9D�Rw/�?j��̗mK�;dNIy��&��a�ٽ,o=��	�$14)���I؃��aR�[tǈ��|%lU������"�&�䴠:������}�[�C)�d�xf��ܲ�y4c�H�j
���d���4{���b�Hkl�M=@L� ��|�*k���tBy#�
���C5d�UG����V ��>�Jn%R���UoQ��	���٦��ސ7u�|���9�ڋ�7i���N)��D����i7C�0��T�f�'�͈Xn-'6���;�cد��SC!҇�!� ��l���EN�cX�:�_�&D�(����b�t���{E�ߑ���r;�eE��auwи���W{s:��ڝ�bd�Ŭ|�A6�.RW�M4�$q���Y�g�G0L�u1��.G&"⇓/r4���3ع̮��f�(XlxVHYEB    4089     e40	���:�:�ֹܲ>���sNx����Y �P��G��T�v����7&����q�D��vʖ)V<+�p��
w &���}\��O�!GOМJ�Ab����9&�y���QLq]�@�3ϳu}Y�Z��zeF�q��ا�ҟ�}4�3�Є�f�ŭ/I\��5�2���ky��G;6K{�e��E�A��JYJ���C�e����B(�Q�0k�<<�	�
��,ՙM�����#=<�M��y!�n)�ki��	a����\�X�9C������My������R�J �(��Tc۸X�|��(y,���>�J˻
^���W��������_�J��d��:�;y��F����cw��+���+��S|F�P�˭�Q��ļ����4o�ފĺBńs��\،�f�">�-<O|�{m�f	�Y���N�狎g���W��b*W���:�Z��ҫbm+a��io�}��k�	}Z�ȹN�����6;ǩ����~>V;5��Z׊��6��3�g�G�Byr��|#�fap�OX�rv�S'���� j�� U���ɿ4~����iw瞞V�u4 
0m�n��.���Db7��@\8H�Cp��aȘ���ż#��tVO�3 �ECTA�C3k�.U�r�HT�` ��^�.3Z��m�3ST��>�#dD�t
;��]|�f*�\0��P5I<m�(.l���K��IKjA-ȶ�D�,
۩�3�ß�o�u ��J�Yáp��|L��6�x8b)�$*�Ǔa�
���*B�u��F�*��߻?�ǥxN!5�Y� �J�R���2�&�굥�6�U5�����V��J�nqG�K�s��n1�[mp2Y��x��*t���N���D�fl�_e5����I).Ӹ$��N<��/�Sծl���{��w4�If��'�b�b�M_Z��@g�Fi*��9��92���%Q����o3�3W(3l_��>��zq
ќd1mq����'P>.׹�(d��b��X�Q�$�
��װ\��7���T��&+F�5x/���p�@=�N�q�������?B �А}�H'`���]�t_�#7�(n�2�%������^���f!��j�4�|i�w2� *np��r� ž��Z>c����y���٧!�W�H/���E�mX�2�]٠(��w{b,-���-u~%�c4K̻y�~A�~��1���9x<7���}����A������N+炷,�3n�����J�2i�O�
.�B���6w������*�ԌZK�{�A�Ū����V�z�+.�����Ǚ򑦧㠂M�hDx	�<���
@��4�WWૺ�~*V�AH�� Ԑ�q�
L�
/��9�֪��M��Q��\��p����a��wS�5�c$lK�X��I����Y։�ዴ:r+q"�Yܭ���l�ͨ(mq�b�����)Ұg�tQ�֞bC�hX�'"b2��T_��e����i�	3��0�-�j��h��+�ڃ^����:��D���[,�L��!�lAQ�ӕYT}��u�I7�}
Г{�?�	=��a��8�0x��Q�f�W�3~�Ƅ��Č�\m�r9��Kz�q�J?�Sm[�[~7�= v�K��b7��]<5j��-�.��_S�T�}E��mi�a�d�K��JW�r�n�bI�%�M�t,�����Lm�!��A�?���#�+��Ab�����K���:L})˻$56Sa��ڊ��`ă����(�1t,n���~��T9���y�c�/�`��s�XfC���0G��P,��t����;1�a���� ��Ʋza�@_�j��7ڂP��dtr���^�*�-�}�q��f���Ҏs`��=C��-���w���COs�7yVc���b��*��3\���[�\�D,ƛ*A@�.B&�p`�\!�2��]6�G����������e�k���n�5���o��'���X��#$<N�Ƒ��̐�V���%v�Kt���m���2�|�$#I�����	Eħ��(v�f��iX��w#��*񁢤������%�4�����������S����r
�aj(�њ��Y��Gd������r]�Pp�&�9��Ci�����s$$uG��m��M�؏���ß�!	��5B�.!�n�	��4���	��'�����q�3UAd��:^�����&D�2���l�VGn�C|-NJvHF��Mݔ��p�F�IQ7���L�^���z�D���!V.ۀ��2�ɫ��׆k��>�קQe�Q�g����w�%=J�W�;��?��iߞE������k��A����<�K>r��Ql��%b�������%��_w)I��x�r�>�C��� ��H�0�W�甯�c�Q��� �~��*a3N�r0�1l|�]�=&�b�#U�[�
㇅�n;���|�,5�uB7�"���[�����c���р�����G�%��ڒ_��� ��5�&�����T���w��9�:G�pW�9��Q��}>��[;[�^�3G�����%m�lBLi�g����J�Х`����z�_c��O�r��o�?��u�����O��ͬ��	˼e؆���R��oKI� ��[P�y=��O�ڒn��L�K��ی���㽩h���sw�O���(U-�H��9��եMQ�.�Jq�R���Y���`Ky��		�� %���� �8��^+%U�1����ĥ�4�UE��C��>�_!/wd���tr՝�z`�����Д�X���Z��D�d��9ʼ��n����J�RǇ�nW�Y��;���֌ f���ü1CP!vi���� �L�5I����8@�W�#��N�Q�:%��e�-�N��*�k^=]��Q��}ncu@��MoV��lp�5�C��5U�����,�ں�ٻ�YeƑ���*G��f��j�[��ckm?�� <&_�z}�L'i7�0����3�-�ï�C�Wdxر�}���Tq�t�&M����W��B;��Ǽ��>$�AP|����KG+����nJ@� :��6k���k���}g��G��!>,��e_4����c���tjGD��- m�eMC�~Z�O�V{�2�jk���$��"	T��F5
�	TD�n�~� �"�|���mX��eQj�����A�q��O.�_r�@����ך�ߞ�=���ΩY#-Ռ\M�W�8�_�ot$�Y������m>xP�?`~e}�����Ad�ǆ��>և�9��0�R�<ܹ� a �^���Z�_�0�$"`x�X�b6�R]:"yB%k�q��Q`6�����%ВvJ��"Xb�h�?шhSp=���^�N)r���e��C�v�]��$��-M���n��� ?^R)�id���W��#R�����Q׽��<�!_\����df����,�cJ8�IW����.x^4y������YS����ESK�ׇ�α	^`�=��wR���9A�(`K�-�X�/��ఉ����6����uc���C��Thf<���$S�;�t��������I	�	�j�W�+x"�;�d�2�4�GN)�~bs&��(a�yJ?��*��$�"˚[Xe*b��=T�02��d����:���뎆���hY`�