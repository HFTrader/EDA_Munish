XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kɸ��u�4E^I＿i�"OF w+?-[h6�����+�+��G�'T{;8�7�4�*�-�Z,�����kP(��qP�^��o��'*�{	�J�_����2�Pw�p�s��
�W�6�eo�!%��O�ь��8sq]6��g�ڎB"}��ǹ9j2����>�o�(�G��Cն��ҏ�s�ܧ�}ȧ�c�_�x^(�u�na6J��,rJbĞՖ���8p�-W�r4ڿ��I+=8�?�_��D5?.�F�6V��.['�����]�H4��Hc\��
�|:m�
�E{�L&�k�1����1�~4'�/��."Jc�%��M�JT6�z�G���!c˂��5�F��ʴ�����|�0̐��}�Oa���ϯ߀���E�;�����9��`ÿ�~W�H8�t	�.60ߙ�3�B��׬�CJ��o�;<�oO�̏��E�;�Uq�8��y�3ӓ8`3�������mU�1O`��a#E�#k�����h%��.n=���aĖDұ�7�lkey0S��ឞU�.�m�}���z$6󉥘z1�~Ċ�&�@����]�C)s�a�w����"���c��`�YC;.M�wO]m�A5�Y^y�?���:9�N��gs}ذ)w)�"T�Z^K_��mt�F?���i���f���֖��Vp�~4���U�F�o���Vi|�&].�9xrZ�'�L:���1�6��fS��l�3�rh��R3y�=O�J��h�F!�]V��!Ax�y��x�%Ö�XlxVHYEB    4052    10f0�%�q��8s��d�QbSru��"��9�T
���g���M	�}��+�(��ZF�SA�_)�aY�W���<�����S <�s'����7�k��7���ۣ�����9���USFX���棯��D�O"~�{��d�LCn?�d�X=�+I�7�M,e�J�Bo�F���)��v��K�C�,��_C�5r�Yj�����GPE$�S�^����樤�2��z�"����OB���U�l܌�ON³kNB@�Ŕl��j0�?��5��
��F�`�L��V�yU!7N�:���k'�����@P�&����k5�*5W�#,�뒶��VDg�ęb���/��85Z+q-��|.U�(X^�nT5�Tr�}��3徟IAX}y[+'W�"�!
��E���G��
6nd����wV���1j��M��~O��]X�yLRokv�.�0�oչ�+�������)�L���@�{�XV$�ZE��@.�q�������+�̡�0	+�,��se�(D��<}���kT6�̎j)��_���5������S������B}��F2"�t<y=�ə�;��!�8�GV����x���5�7�m�@<���fs��\U�)LM�0�	�8v���2�kP'l:�|m��:˃d�g\A��w�/<�{���U��>.�HC.4ʯ�����E�G�������?#V`Z��k-0��Jf��	W�#����Q�ȥ�������x�c�d�5�� �iFm���@W��� F����h�=҄���Y�pQR�'�Q�
����?ݿ�S,4��A��)�5�s����z��eQ��)ˑJ��)���jN�o��3 �r��,���p��v^�#�K9��I�j_,���7 ����1�5��{�{�H1_7�+ў`e~9���:^���<�;k��mf{�g%�`�#;̻K��d�F���K�� `�-��C���2�l9��Gs
t���T���2����6v(��w�Ūˮ�q!���D�����]����v��ҭ�!�_Թ�X�Y��}�O䨛�J���{S�GXv�j�#�hč�1X�f����Ѯ�Fr#(p#�������=u�ԾV	�Mt��v��TCk2�^��kВ�� �h �pR��d�����-J-N W?�Y>Ύ��*!�V����hS�텓���C�%���NqS��"1����;c;V�WȌ��5a1���<#����F� �G�>�]t�c��I�}����^ f���1G6�2E���4�؟�(�K]x�k�k��x�ogp��s�T�)�]�` ����!�/R��@��#�$���!�㛝�h�f�F_�*aw��샌,|�{'�)L��C��7�oQ�qVf+_T�2�Ne|�|an�h�o��<�xJ����I�ZJ���ڄ�XP'�T�s��=�L�8��MZ>a��vy��"������@��vL��G����$��
���f�J����m����҂S�#���K���՟�`M@l�D4ikō��,=Ʒ�;�x��9]�kN��u|���68�;=�խ
Ƿ�j�b�G,��X�>��OS_\��m�v�I.8mD��#�
�W	�� ��LIR�s��V�p^+(:�|�������Q+ϲ:�zM%v��8��o)�:�QU�R�Hy?| �R��Im�\�RY8�^���p��1̕~-���� �]����nw[W�Ȫ�,�H�X�o��_���S�R�^b� �@сt�Dް��.��؁��O�kZ&��ʊ0�n��	٩B1���)d^���E:�,��	>9��3����rR��c:�1dt.��.4���?@�^G:s�A
@�fl���l5h�� q����q�Z�ч)�z�`t� >3C�)Ī���ӵt���iL��|;	Rl�O�����Ұ��e����	�t�ѫ}w��8m�C�s�h(ʔ�����K=��}�A����VW��=��˙�쿌d+�?ui�W&�t��`}�V��m�Ě!�ө{?@��=բ
{i�$&<=��m�i�,L�IOg�z@�A��G��ͳ�[{sL��?��ϑ�C*@%m10�.C'�\R~����W�3r���0)63�s�K�pi�O����?؜n������}��jg%�7?�,��4�q�I���rk�O�7�q�M����W��E�쎔�dh�.��O�%nOx��s+��(� E���Ǹ}T��vo�n�`���C�t��<�@���<Y�ғyDQuU[����/O8���$[d�u�{:�Q`�a�.@>X�U��H���I�~���k��T���Z�u�<+g�itNd�ďm*Tc�Ht� �X���o1U�����k[/k͢��Ӥ��$��N?c��;���Z�呴%�ʧ��PZ,�3���ϕ^��=���W~@��W��Wؼ��`�Sc��%�F6r삻��r$82���iiը�+�z��H���d�H�q4~��{�I5̭����qHY�}��:ArmO}�7�n��2�T	|C�t�X��MB��%��@�$�l����q	�����M$����4�3���W��x�#�Ro�	i� 쩫�j�t���R���LÝ�S��+eۂ������|����|Lʴb䚷P�O���h]�D3ّ�'��.�]�d׵��<i%9i�4���a�~�-�Jߍ�Ik;�5��l�d)&��	�o^�乇���1��iB55���MZp�I�[����KJvbQƺt$�?^m�iMzlm��Ȗ>���K��I�\Su�!C7Lҥ��t$,���D� RЕJG���ʼ��b~��-*�Q/��Ʈ�p�ed�m�Wj�X�U$�q����9���MqF@���7�w�w0����Q=�!ϔ&��ߧ+�i0b�dۣ��U ��HA4�d$�7s��f�뵕��a�R�U��8?��ME�lZ���j�WS�<u����-y��Q�2k�r��Cf�Ff�hB�|28jD�q8nI]hS������~%H-���b�s�7��垿z���cj�f��ƽ&�T3o���.����'8�Z�0"w���{��!��u8��q͚ųF�>�C1kV7��2ǽb�v�d�F�.lo�M��2ر��]]����C��-�3�X�"�4ż�0%f��L>��Dtl���Bu��D�N�%��KD��O��Q\l�I�%%�8�����p��1OW������B��\1��I���Ƽ�q�������>u��6u���i~J@�>���h��c��7�I���iK�I!����B5��%��b1���N%i��a��V��K�2����L�F�ӶTi�/��J+%�B��Ђ���ҐS�w��H-�y����:a!�r�s�4?�Ny�]?���ژ�0��P0�tv�P[�������BK������i�\��P��h�[�e��Yro�e��f�mP2m~2�����N���=�F�W_�~�� �7�	`* �|)��[�>q+���r �(�l@!�/؀�eW !!oP����eF�mm�'=���B���a�C`��2�a�`̧b�D#���c����pW��%�<�� *P��r�(#�D���u� ��>%	��ө�)z��:.40#YL��fΟ~�`�f�V,����RȂ�`�+��1^��202�"1��?V����P����!�Jq�sP�Y�9��m�ǈ��	��Ֆ����(b\�05�m�4��������*YK�h��wZ�c'�T� ?7w���2�ݓ1T��dj�/�
��f�hzo���h����&5�&
���i��w�/��ο���Ӝt;\��$v����ͮ���Dm�p�xf1Ɩ�Gg����n�[���vBC%ħ���(��u��Ŀv0�U��5mr]E5�xE޴�{P�1~�����h��2��~��A.h�2
�Ke��<�H�{^B�&M�y��Cr�l�DdʬB&�Z��#��ͻ�Bepe<�T=P���)��e�-��9u_��2��{���DOW�t�#�2o��1�;���D�b>��N�^x(탬��(pEj��c��_���p��r��==�&z�܏��0���q&d�quG7�b����w�/D��R�>s� '�đl��,;��;(�<U[D�o&ߥS	.9�qSņ_�԰��7��{�9��75M���_��}iM�27~�@��ۡYEPma�:%:�4��1�
�Y�L�R����������8�ԁ����t����ûxI�?���7����o [-�w�8���