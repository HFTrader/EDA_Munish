XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Eh#M����:����4�6��	|�d����<�o�N��}���F%��G�Zp�������v�t�ǒ�Yz�8���_=����ȿ�j���9HD}��,P�C>R+l�`�m��*�t��=�F�� l��$Vv��f�1��㵧&��ܙ���f�T�X��*��Ӣ��\�m�͙Ɏ��đ9Ϻ)�Uj��l����S�L�n"(����53_�'��A����y�SF��&*�ب�������u?4���~��e�P7����z��G��p�w0hҖ.��r���J.�]��ke4��	�wӒO��3p���	��>ZVo���%�lm��:�Ǜ��鎖O#�^vw�[h��N��P�/�m�2:U<��r�Bǣ�x�0y{���M�(+t�M�I&�)!bEz�g��(<!{��L0�A�����ҏ!8m�qL���&S3�Fr{��}i`�i*���Y���~��x�I��u(>��|����Ӟ������rf�)���dq��	����n��:��<8 ���ަi������u� x��檢J��ß�E�`G�4B5�j�	�V����@�;���A��KA��'��<��{���.|ۣ_$�g=��=����`��J|�Z�ì J�)�ƨ����[����	69���aG��y5�dԲ�é/��]w+df&�xj����KtBT�}�d��9AA�����J$xjrZ� 
˷�.��`�ɽ^Y�F������pK�7Sň_�ɴ�^�Q�������L/�XlxVHYEB    50f8    1010~ߓ���&cx���R�u�Y�K�\d���L�G�\5�> � ��I^k�~�z�Mӆ&���Te�Xmg_H�����uArt�<�����lК!����pQ�_�.S����>k%2�Y��2c<n�d&*�?>]�4 O^�<$oм�K�Y+�c�Qĭ��4*{��FͰ�a�f�KRG�J�=c���{w�
Qo��#!���@G�T��k�F��1��/�/-_�T�B���,ذ"��3p�������R[KV� �x/��X�B��\5c]{ؿ*�A����w0��۱:���6[x�(R8i@*X���j��}Z�t�4��n@m ��8�Œuh����>�k�����gS�epqY��7;5��7��8A]zϔ^���T%FY^AZ��gś�AfJ-ʎ��.�k�}���^��� �9}A���S������Շ�3� ݘ)���e��>�]B�{7�YVt��Kʱ����GDsq��;v�R����J��y�-MX'�R�l.�z�#� *'�qB[���Z&�d�@d�ó5�.��y  ���1������mKmb�pf�O�w�b�Y��wR��J��:yZY��<�JK?T�	|���������uc�
b
��!s��a�]8��;y�V�O��^����ﲾ}��ĥ���=~o"cl�RQ\Ĵ{�%
o�)v��Śi�Z������/�U�O�6�K�P�u���}E,�~de�h�9��b?N��/����aA�w@��V�������I����x�0ۊ��o;�3�JAmҒ~�8�t7�_�Sg�����g�~]��y1��@�a��Ov����:y�=T{�|���,�{�p�򈱍����1�l+��g<��'.~S�����h)a�z��uPߒ�-�X�o�m�(��)���Q2�C%��TrJ� ����n��5�Ǭɿ!��i����+IUM��[�Zǜh��9�@�wA�\�?����u�n��kv�Jt�_.3�v�M}:�j�1��e~8`�_Glq�4�*ZK|3߰��G����i��v;+���>�,@<wh`}�W]���W�]Y�͡��uY����^$�}7�L]��9!ۢ�s4�d�����J[Z�j��x�Q�`� �Ɉc��,�y�zf��J	�GЙp㺂���]�ƿk�߮T��^��-3�0�����z���»NPpV:�A5e�R����,����Һ���+S�*=R�щR��|��v�9�.�b�����\��pJ�pZ@Pxn�D	}�f�����8�z����q�!�:���E)���7���)w������g�Q����)Sцf71�檄;cI���P�ؼ�`�^�����
$10 �C[�_CKY�'[�|�^��+�q�;@�����i��,�\�1���_ߍ���*���'�P�*{tm��g�y��M�_��̰�DwC��d�ptkh�ck�A���*?����a�X�\�5{�������1��g��.��C���Sޒ�ބ��![��%=�v�ZB���xe<Ơ ���0}c`�^�Y6~��A��� 5�L�!�)��)��/�*��`�ZQ�����9X�MD)���\��y�͢*"D?b�����=p-�A�̍t�,A ��� E  Ft��M?8Q�wa+&�w0�N����v�z���7.�;���e���?,��>���k6>f��*'��j�h���c������ ����,�>\����9�=zQy���|:	t���j�O�3xDJ�-[��������̚���#&�\D�i;����Q�vD�v�n�t�nK#�c���ZU��27) A˗�a!�%jI�<`�"���[�@33�@�eHzNgQ�A��\���Ĥ���θ�$v>k�'��`0�bʊ�z=�ʅn��Nlb��|��
�~����`%��y�#{��d�!��:\U���=ߒ�T:��d�:9!��:)̦��n3�x�3`�#]��,���f��@��V<(Ŵ8`-���e��U��>~o��~ºo�qTRG
�(�k$����h �H�V��ʂr�SoKu���TA/\���B*�'�x)~/W�4�*tV�(��L��u��dt�	���֦U�(�5Iv۾:n�(�p�J�0ؼ� `Yâ&�qYf���:6��Zb�yzЙ��2>��.����O��Q74���7�_��4b`Ly��Zu��K�;yl ��.U/2S*���|X�mb�w�/&� )�6C;f�!m�:�)�gG�����J�CB�s^��|H��L�UR�HBA�lX��(��Fz%�1��>C����?����Q�Lh�/�)�a�$~��~"m�������O�?�}s�a}���� �w��r*W떊=�$v-x9�c"��֕ᬱl3iN�T����Nw�Q��2q�ܑ��s���Ք��4������i���yS2_�ح	�	�5FF�X�X*z��DT�_�IZI	��	� �SO_�C<-��t��e[/���%�[�dA��/�t��j�
D.��|1J(�4vٖs>΁���]ܨHr���J�s��Yם�;):�����\��w'_G��ԞZ�@�*��fK�Ia�,	~�y�Ĩ���#���e��P�`&� �µa�U�)&e1j���~M��%Be�s�@���jݭt�'n@��=q�X^�yͮ�E�+5�;��2>f�Hta�fesQԕ���!��D���1�j�T�%�Oc�e����Y���)�9E�ls���:2nH~�&3��� ��H�&�*_��(|t�	(Bn(�DTB�d�O:�G6�\4C��.�6d�}HJ�"�b�]c9w��cM^M�����Pf�q���v(i�G���n�mv���sA��;K���Ss���#�	%Q:���*pf:\�m]��3��[$çک[��:l� ���s��o,?&���w6��CʸK�4���?|���@��W:v;mJ��+��{��\�`�8#���J)��S9;CF�F)��3>l&$��o;��VD��e�b>�n��ⶳ2��@5���5�`���v:����"駧K)|p_!.שV���O�;Ò����])�q��M�:����m1h7��\��$W�8���;�i�DEڊS\�@ʬ� �
����0�����V���P7�T0���C�[x�2r���;���W�:i�����3��(�_�2�g���b����<��r}c�7<�36ܰ�&ؘ����M�K7��+���Qݯ��ʿۇ��u\��L��]���F��|w��Y�Hpm�a��XvO(С̨-]4D�͑Q_ޔ�ܶ����7S}�Qϓ+�g޴|s���<93w�8�'�#65c"��G��QcNٷ������| �����"�ٓ#�o9��.�Q�%��RO����`#���4ozC��۞Jt�I�p�G�B�YF�x�~���������$�o���b�$��]> 'd�Þ�s$�_v��UP��HƔ�?�㚋��e��]�=Z>��ؕ�1G,A �B�ʦ�Y
�s��Ke�?8܅�"��*�U��Z��$u��.�D�o�����:f�1�)q�s�iQo�Q�R.ϹJ��TG�f-�>.aMF��P����z��7kp��`cr�@��y��GI Q��l��/Em.����u�����)�,6˰�Ɔ�R�	��>�����c-�p�聊֢��k�IKD�(�dS*Z��������\S��c���x$�1��L�DO/�Zb<�*�2z��h�� }%:� N�[�c�hG�|m�D����Z#E9D_Y"�n�����2U�®ɴ�� 6X�=�Z����	N�h;�%8g��z��:9�����a�y̹e��<��K@�35ak����[��[���d��v��1Ǉ
8d6���-�k�78�"��a�.�9���@^��Q,|9�ə��:���`8��۴�;���H�u!S	f�Ϭ:�j�Qٱ����&��,�iĶ!�' ��c�5l� �l��3��WEx��<(ر��+