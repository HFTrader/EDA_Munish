XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��LDrŗt�K%�J���>��b�,�q����Ax��GUdw�IW�q�>����W���[��5�ՖB�(��]=�)��ރm��w�ނG�IG��m>	�R�n*ǹ�����Q��r{άwB���������n�J7�9�e��r�9�c\�d)'��1)^��%kZ�I1k4��pF�C���&ܬWb�^s��Q$,���1d ��^\�s%d�ԟ��I�{f����4��ڱX�=�r�%��\��W1f�6�$-%��Ǽ���} �ӗ=!�+�ꀥ��ƕ�-�%͓%�j`:V��p�Д�j��Y����6D#92����;����Z�-vQ�����K�݁�Z���6AW~Q6<G� ���s_=!6� ��v��8�~��_\c�ꪅ�&��^M�N�a�Xm0�T�-�}��N�	��c�	~kO�(_����y�~�A����GD�q�e�׷��~"�[S���`�T���׿0$���3>7�D��i��6 ?GG.ɖ��#V��n�4 �?@�K��sm�m���nr���8�T���5g���8��_�
%�Y��i=��23>l�1C����q���Tgc�7��B`_�d���V-���(���Q9���2�n@�'���==
v��2���#���.��eo�T~�u������^�.�&���9 ����;3;G.M���MH��K�	\Xv�:qAl�#����g����C�ҔZ���l�lE�
���8%���J�l��~S�XlxVHYEB    1c45     950�0wr�C���C_$�V��w��2Kj�J�r�[�Ze��4-4�E�U��a�N�٪3�Aݕ��a��dGf<���*t��ȩ��6g��v&u}��֏��8�b�aͮy�n��rk����RNj����9�T��v陔u��O�Re%o8wQ����p�Y%��R��U�_0z%�M�	M�Dh㏌M��'Ms��y����<9��;���k�<��/lǦ���#����[2ퟌ��b�@F����Qg!g*�c4�	�w��)��D��s*^C͜�����������S�,����{6���-g�=K����<���"��n!q�ɛ�!�d��@?�5le]�>j���.?|�wУ.+�K�����������>�ޟ���1Đ��#��Z�C�kg����[��Ѵ�R��N{yeY��c��%XCE�He�[�{�x���K������҉��g2�k-��� �dOt��6v�� �OFTcd:�#��v����2�0����v��b�4��	ڴ"����\-Bj�9���V������t=:;���n%E�����'�#�/��į/8m�?mx�X6?a�a�SlR�:�~iB?ɃJ���ס�� ����T�4(وDzF�u��_Z���o]�x'�Q��V�`hlY�X*F)�d?R�PG��w,�;X���,�����hp�L�����k�ۛ-�9w�s��P�~��A��tH$ ���g�]�d��M>�%�!�^;8��G�Jx�]<���B����@��O�-~7؆*
� y���5
�z���xwx���_]��&���Q�s�T�b�1Y�יu��|��^Ʉ?r����x��$���ύ�O,��?CEwdg��Y��Ө�f��z��cfM]���V�����Q�^��#��;<����*Mm���\�d ���( �X`�7P�ʒ�曙d6�8a��ƭ0ҔB�`��*�Ӻ)Z|q ㊽0�f�دʇVӁ��~�� ��{����� ��� �W��Fo��K�׼Ք�>���.F� �+1V%�0������q�91f�[���b\O��ޟ��Ҫ�i��m�T1���Q�T9��(���� M����.#ap>-�zCI*�dQƿZ�Cl� ��ae�H��B����1]��2<K��8�oq�HG"��}��G3��n�eP������h>L5��9���ahi��,@�6���R>��� 2���X��f�d_$	�B�)��Jӑ1Y���v���3y^d�36��+s��!�@�R�[�@z�Z��8M2�s9E��G� {��I��Ys#$8ą:�M�j�˨��R�_-��a��BXP��<9�='Ž�J�N�Ǫ�;����&�ϺP~K3{?4��1�5>+�`�g���)�L� 3�C��S���� &�cE��m�.p��_��7=��y����v��3�-K��͇l �$nWxc����coG;�ǣ�|O�X��v�t��;�V
w��%�������$|�Fv��I)�_�k#s5�x�A���aZ:i"$�����]AhLZ��@7N`:���\�R��|Hm�Qҍ�V_�rn��K��sBF�R�{�ȄI�ݟ�i�e�g�V_���'����{t鞋�"����I�t>?jX��n<�ƞ"�����L����8�G'�F�uY�$�~��P��n85ib����է�$�ˎ��䶄�#�<�=X��� ��_h�-.��"������*rC��k0���zTS*�&�_t�$n1 "��U^�aĶ.C;�o�X�ԇ�F�d���u�F��;O���>bl�qK=��k��5�w־�wG�Ym�p�P�@f$4�2���7�8�~f�u�B��.����-z�G��Ҏ��L<LY��ٸ�x �{��r4�{d�OЊ+���W�D�ݹ���)ܟe���[ �����:�Yu�������l-=��etEX��a=[�~�k��:���F�5��I�v��;j7�O����ddk��� ��
 ��i�e�d�}��w�F��+���v�'�sJ�Ul�,CRǗsVjcoO����I�96.B�v��Tu�U��oH~hU+�w'v���;ѕ"W��&��U*��Ko����V�y��D�p�����`Z�RO��UK���HK7�����u��bL���AcϚ㯋R����#1J��O�x���m2�����!�{=�EL��uؖ\.��b���\��GC� 	\2RG�S	��X�hE��"�� �"����&�dd�\F���,<�3�ខ�H{5F�����CX[�:& �� �o:������BGh8L2@���)v촖r]Bbj^��dU)���u�