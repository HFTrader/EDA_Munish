XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��+h#�v4Q����v���g<t8�n"Gu2�ߐ2.lχC���*>u�GJM"!�Ҏ=�߅��h�*�ǁ����ys?}eUZ�L� �,��H�Ӱ.��z
1���Y������,0�E�8;�����K=hq������:h}�`�b�(lV���y�Fڕ*��k2Q�aQ��v$`�ì��ńA��y��t4���NJ�hx v<���`W_�W�yֵ�i�\��γ��ims�ir�4ܹ���9CQuxT���6�3�r��OR�Ys�,�i�Ro����;��4	.�XI~;Q O�Lg`��H�FNt�H��W�3/����>����*D��o���Le��s}���/�r_�9��lrfvMf�\=$dKq����a�O\]�ޫ��$�|�B� �.oH~����uCu�6ʘ'��>ܪ�T ��3�#rh.g<.0��^�8��+��f q�W$v#F��}U��l�K�l#�E#I�A��-R;|L5�j�0:�I�c�k���U�i0WS�%���fyI���u; �����Vh�s���X�1	���f�:<�Y��ۣ3��� �AL����:K4������g{ٟ {���.Y��W��k#�,W��i�@�=���"U��8��Z1碅4I��Xo��V�>ީ������#�S:�5ۍ�8��rQ6� ���_S��j[D��S�0>��M�D��]�U@Kjq��(��ɥB&����D"���q�C���?�=��u������ྩp��[�����XlxVHYEB    9193    1ed0���q�7*JB#��@�/f\�3t��=u�$����VF��G4��|�^����c#��75��w��kGS5�@en�	{��e�H��*^��<��(�{�Zn��?[=ޛO茨{I2jR�����Gӣ�}ڭYB�+*kٺw*��>R�ZC6��)��2��
N�-�<��[\m��L��z�,D��y9R�sGA%��#]�AkKN����RϮ;��i���A�7v�eDf���l�K�☨�JM�x�I���f b�/r뚶Q['��/�{ǜ�-��FUi���bj����L�;{u��ͮ����T����,x����|�!"d�%�@�G9���ɔ$D�M�+
N�19���w2❳NW�44�ɔ����W0��|�q����h��?��.N�e [����}����K��$I�����J.!"��� �²�.�W�����\�#E���rt���@ܡ�
��8�I/�ag"i���d�|Ҷ��}�ґ�KsM$��(�oK���i�ٟ��"*��x�ǥ�&��ډ�o�!��ىN����9po��UG !��Ս5H�R�h��39����[��E��Q~Ҫ&bVFd-vZÃ��O0�8�fG�.��ڙe�,]��/%��f��6W+��q,7�Μ��:��4�v�)�n��)R$�~�9�_HT�𲲊�b�ɁO�k�0�mǼ�I*�={���#��g�;�La-�M�B9���w,m-��t-�a�EI��\�a���j2�·s���O�Uc�����/�!릳?����)�VM� ��l������x�v�b�(�*�E�؍^@P�\�2A�A��*�_-6��R����۴�\��i�2�l�TI~޲uA�&G�<]�<>!� ſ�9J��>c�n��;�љO�q��� ,�x?ЉZEyGc=����iGfF�c�"澢ݧ��t�%�W������_j�Q`ŵS�=��L����ٵG{��j�����\���u��=e����u����s��= �a*�u�;J�ڈ��ߥq [�G���)Gu»G���jgmfP"�	ĝD�4
���EΑ~�)�H���Y�������%^b�i��]������eh�H*U���s��cE�gR�K����?C���1�{����2�mљo��!SZ��Re�ݳ���B�,�����뫩2צ��T�f+ K�!�����t�:�`�=PƶW��3<4�u�C��s�8$Qv���Me8{/Mh�ѽi����vU�9�!�5��" �l�I��R�n,W_���tl�\*�X�<)�.�YTE�eF�ͨ9�kv��9��lX�௡N�B��G��*�P����϶Ք�.`&�LS�i�����'C4A�@'�#oi�y>u���̙4;���Q'���˛�����B���˦��gw ��kl�dʵ����n��C��,�_�SlE݋(*�W��q�^^)Xa��wv�Rv#���3`	�n�M�P|�, ��c��WG�a:s�?��Q*<���*u�9c}�o�Q����I������W���ۨ���vpIݒ��/ĺ�V���s��b	�t�t1�Ĳ=��&c]ҩw�u�=BZ+He�LW�:%�~p��������6��sl�9�ű҆�Dӡ6\�Xwoqw�X�7��c�Ӈ�b|x�s���S?;L�U�wK��.X"�nnw�o�W9���2���P�&p��U7ib��1���?PU�� �Ot����c`�xF�	NW9k�7�\!ȑ�O��ҩ�tq�M�	$Y�	B;*A-��qӍ|�]L�G��O�i����N�F=�׀cQ.׉��c~p6ґ�� ��d2���{n�S�e�O��͐Q�}H�^9#�!�HH�V���Q;�J#3���l���L �2N���,��'���i����T|Dm�,l�0�&�'p��71��¬�.��.���}V%���/@�\Q6��q��D����yxh����ZCC�86Ӆ�w�7��*vzU���
R� }�
J��	՘���Y��^}����'}��bu(��D��wp��R%�������M͜��{��Q'ɂݦ,�����W;�0+!Z��yI����X�x�D�/�>¶�طc����2?�d��B�`��9 �^ȳ�=w zq�V���*�P�ۿh����.4�g�%t����?�<��1��+@\�n��k<���L� `1c�3%LLdEK4F`����
��B��:u���p9F2S�{�K� �hw�e��.-) ��e?�Z��)f�J$���X�z�v �s�1@�Gp,��	��>#����>d�9u&@��@k+�b&πl�l�a7����3�)���0� L�`� D���[��_#cU1�7��ܿ4�z�מ^U�ѧ�q�.��C&�N��,sJ]i��Z_W��ht�(�O������e�[��^Ƭ�U�ME4�kӲ������:D4�\w)���B��"ǒ�$N��.w)
��=�Dv�S��d�O��3��DNw��?�Ӊ=��B_�Гr��3������?����p|G�~���?@���<�-?'[u&,tGr��%Uja�1��{��N`�*�I��h����BLӥ���+�p�UX������5 /Q;�j�g���N��Os�@����Q��
�����2�
t�p�y��;?iw�t+c�J�)<)f]8V����^��7qC�_��!�8ͥGDu۸5"���,��#�h�d�\v�dc�ջ0�xx�N��%
���MMf�s��r�%��_F>`�j�s�6:�a��W\�<��n�Rf�6��ۉ�aCO0�E"���*E6`6gm6�NJ�d]F�V��3���O��%��ބ���	���AT��ݝ�5Z7����9�l��.��		D���r�������K��Y�E�o�|�ϘG�?CO�bW��`�,A�O�~б�Q0~#eo�rO�=�	�8�����5��JY�t��	��*��>ȋ窮 ���5��	��W^���BX�w�D�"c\�X�E�5�"l�����Сu �:��M��Ϸ�[s���H92Ck�>�"��D�P�_�^��
��fь ��b����=�d����^d�����j���+�Z�4��>>$9��P�U9���B��d��Ie[��;�mK�=����j�p���8;��C�����\�D<�uM�U�`{F,����yq~	":����,�V�U�I���
�P�X��%�3�!��JX$_�@�*�H��A%��4B/K=�2ÿ!Gh�1��a�G�S���s�)�\�a�.�;�ځ�:L@�K�w�����W�>�F�JWȖ����P����Z	$����Xa�p H>Hs��[[�u�ep���P~�:���щ	��0��+g+F��r�x�U�F��C�J�Ѝ���Ͳ�ʷ�I�E�����_���'<����kS��(�Dxok�!�
 R�sj��"��a�F,�*�������^�I���PqW�Cp ���]0ٵA�n?����uA�Bֳ��3ЖH�:� �ۮ-�y�k��˛�y�e��s�m�v�M��#�st� U��I�ug�!y�;�)o)^��rU��2]�'#B�(�N.D��Օ�ǈ�����k��G
�ӽ6��PI�u�-܁��{��9�	n���4�9�H��;6C�^ȴ��qW&�q?�X20�[�A�.^w8h/��&*��.����������I�Cs[5�-	���>Wy�P4����i�B�j��ɏ�.	�3���Oa99�6��C1���&��"�A6
'n~q���\퓵u=k]Y]p(nCá�R�Z9�W?�`�'�f(ϑ?�wH�G�.p`s�I����Rن�塖��X��iO�c\��iJ2��6Q��[�[�����B�Aw�y����Z�%�����H���y
�l�?���_<�f�p�n��i�Ru�OJp���ȵ!y�L(.�K��8�iҁQ�j��s�+�%N��ҹ��tBzt��þ}�<��)�IټCL_�;��<:�`��D�ۙ'��2U|�J���� �&X}ߨ���`�~��YHD��A�-�V�@��c���Q�h��Y�K�"�������t,�U����z/t�t�yF,e�f|v]t�)u�xe[(~؊�GJ�N���On���Mľ�3��]�62~׫��3=��m�Yŵ�� ��*��&<9Z���B��}墰V��Ȭ�7���#���4p��y�g�DX$�zJ�6H�3!\@��ܚ�����~H�~(���D��Y|�ϵ�&��� �,�4�v�����V���/��1�f����q芃���e0��<��Ay�(�)�Ŵ������1�<�)G�B��aQ�]jz�Eg�P�����B33�f�����Ź�,�wvt�&l��G�b���ꕠ
�g���R������zG���"�gt�T���0����		����]���0�W�+.��m҈�'��=�s�/��F�y��"H�-#��.�_��o����^C����l ��]��Fǋn&�}�N4�(�_ucE��52�#�������_�q|���/�ivf��EG�)`����`��JT�nʆ���fEQ����"�yOwm
U�17�F�����Mȝ��0�'�J�S�d��qm'- c�Hl��/2�J��YPt�@P	Y\q#x\m��멏O{}T:��(D���,�h���=�:�9�]��M�A4���u���Ҭ��-��;6��$�5��y����ç�Ҷ���m�C.3C�G�(?���|7�t�o
:����J��6������Å��P�N_ߤ�?P�vꩠh�=�Z� �;��.^�DLEe�Q�Q報𵌌
��E�TX�b������_�×.1ϔܱ����ީF���n%����ܕK�Q7e�4���E�ӸG�����P@�$g�����Ozg��8��$�S���k��Ц^��£�/�6Ha�Fh�h��k��᱾xoU�@/�lZ
���T�����=���`����xh�R�'U�N��&�bqz *��t��'�����`�Z����ҠK�6(�Ѳ}�ิ�5��$0�E���&�X6��K�P�6��K�&�g���`J�Z`~2��4�e��ےiq�����ES��S&��Ȗ�]�+ȺǷ�H]�p
�N��)3�����~D�Fy��RЇ�$��������z�X���&;z޿�O�.�G�k���a2��{n��_.�h�-0����z���\�g9*��Um5�l��)�_�yU������t�N��!z�N�ȣ�X�2�´������Jh�5!K�f�e�����z^f���v�������g�zq!��
��6i��1��r��iP��[	�u	A�+i3�J��A����!��+/�qo�3�9�~��@� 蓷xsc���Q�`Ĉ�����=��y� R�a��Q����4me����<�E���#|t�P=��A�WQ��p���!��n��V��v��D�f�$���5/�ܱh -�2�m�p���t��$?�y�h�c<��WG�����+���C`?������%5]f���Ł��un6�dW�iB��,�U�%���t���m�ݰ�&�$���Î�hswh�ˌ���ΰ��uK�Y�d��*�s�(\+}���,�5Ɣ��I#�g}.�s{��݆`�L�1��J��fl�
~:�.���J*n���e]m�M1`6�+v=x	�@���2�ݡn�{C?�K�����M
ck�>���o,���ƈ'p��r|�`_��{�Y�!��D��3LWz��J�����w���g؈A��kҕ��M���/C�H��{���o%9�X��X%�}e�~�Q��޾z�Y��YuN*w����\���d���R���H�pR�M���v��g������N�0Y�p<-U��*��.�5Y�:N��yI$�#�'-�^�xt�9�{�������G�^��"3����mr���)W�����2W���Q���g��Ǝ~~�M��E:V����|��"��&v�SZN�?�:n�$�G�衵�'��tu "��x����=s�<\餹��ܤ~4Rb��D�C	X_=�0w���Xz�Ut(�����Z������fV}��3��J�hʩ�`7�+�ٌ(���a���(:;FX�_��X ��
d#m��9�v�UR��AQ�?д��(h���^Y����'��������8��s�<��!5����C�f7^\��X�_ت2���a^R��3'>��'��d�!��������&7���Nw�D�n��g���
�~���C�[�V�|�W�íF����I��m�! ��3�9@�*�6�b�ϝ�Lx�f�y��a��K�0� u~3�u݅O�$�?=:`��8�=��³w������.��K��U�9Z�N���P i��-;`c�j�.d����� <��#�� �񻻒��`lXC˦?8W[Bލ��߯Y4 y�d���p�d�����$t ��Hc�;�o$�!�R�a�d�T�>�� h��eAH�c/E���U
�= �8X�d5�f֣�Do������+O��(v#�2��ur1�K�ڬo�!���G!sM���$�F�k��[4};�����%��JY�Lσ)7��`4E>��.̚y�w3���$�"=إr�$���=Z?&���)����9�߿"�e�o�Ҍ�i� ��M��C��y}a��*x���Y��=�5ߗwP�&�?�U�Cd+�� ���XoE���R��ğ?ʔ��,���$�Z/�"�RZ3�0�h������?{�y˫F?ڶ�j���.�(J�_�-%'VG��nqE���4�O%Լ3�9"z�O
Zp�.7��Z
�B&�D-��-�z�~���'���\�Yѭ]p7�3��!�G���BM+���ȸ�sm��,�K�XĥS��Q���S�CK��^X�!!���Ӽ�lV!Vg��[��,�V�y9C~���q����>��2��U���9�IR���Ōd���qV���u2C6j�3����5��,���U�]�B�{�-�����4ĭ��4�S�����w��1u���Ǭ	���,��?yF���3B�Y�Q��l�?t��?�⹽���� �y�]�����2���>n��<B#��Q�Bؗ+:�01Rk�k�g�L�����ݿ;ȥ~sU�O�z6�u""h[��$;�Z����=��c&��l�f��� 8�Cx����)���@(�&g�&Q��J�O�n�>�@�딁^Cl�x��ԃ=�ഭ�D7��#;�bx�p����8��S�C}��o��Q�`�k"��Wl��
H:V Ba^?1��2+
���襁��g&��Byk5*Ão(S�*i��1�(�W.y��D��N~��hA����~����$�LI��x�.�6�s�jJr�[���ꄜCVM���7��o�F��%s��DA���"�ZMD��>Om�Chb�MQ}��߃��t�4ZxH8���	��e�V��4�N�!r��ߔVN�j��$��mZ���:��_Φ�2֖�{W��rF���uʇ��XI��	v[�ɓ�
쭬��*i�]��[G7�MA��.�R%� ,	����x�	�=���� %s�%����tN��n{VO�ϱ�D=� ���CI���RЭ�W