XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5���>^wI���v��R��3I	T�g����ă�*�f�6�~�ο-���) ��|�ݏ҃�p�v=�KB�.�E�p~�z�wBM�M+�k���x�-��yCWnӆ�X���-�4�����x��Yg�}%�M�����H�}�ydWSa���3��F� �P����&e}����hq���|:�l�90�郜	iȥ]%����5_{sl���3��������>�������bc�ܞ��-{TU�@o���&v���d�	���~�;�#r
|�L� D}��\<�t�V���j3�����a�/ �sC�x�?�3v���Mо�J�"�q���|�Z�M�k��f�08�V�=����Z�=��;�w��	�!*+��8l�/RL�l�Y����ʵp���S��lb�DbQ�ͽVHq(-e�� ��=Q����K�D׫J�����R�%�:R`�)OKW�~!(�������r'\6�����<�iA�ԡ2m���h�d�bVM��)�g�@F��*�R�"��[�W'h�~7�N�F����A��A�$%�Kg��N� A<f�N<�F�V�-�zo��)�m���z�w�	@?�ػ��܇�o�%kY>Z ��F���N*��@q��?2R?ȍ*[TJ3�u��]Y�q
�ȌS���j�O�����Cw��"	�0/�du0	�=�{�,�jd�l2 ,-�U�Yu�b��Z�.צ�b�p&�'^��D}~.&VG~p�kKŧa���-�u�� o=��&���*B@m��	�G
XlxVHYEB    fa00    20e0�p/V������:��	j^e\�Ja@���]
�7!��RU7H)��*cӜ�!g�i�PC����5�x�srn9�FZ<��X���о(��|GU&���gCB[&��^����?����N�y�f�_S���[�|�d�e��ZZW�"x������U��A�f�ܘ?��!��Q���{F ���uW9b8��wO�&����m�*�!�i^����T�Q(�6�)�:��9�U���-���UE�c��w$2� �j���Qo"��,�Cy��[S��WH�>�%/VS�W�oG�F���8�{�2��vxY�; <74��b��4�f�0�Rx���U�J7�Oj�Xb*8X֞����V52pL��ԅ��D5�*���
1��VSU0�/�|Z�V< $�0���2�-jS� \w\��e�}����j�� �N��5nĄ�&l	��I�(��+ n�S��ۋ�c+(�/6����BF98�~!��	~��^��}�V}�6Z��sAe���� �@�k��Y����E夺X��?ٚ��� ��ю.��r��'�A:��Xy��6$�%�����`������S�6�"\MFN����g$�h�KGֵ���o2��ٛ�D8���*��m{�]�T�I"��?R����d��ݹ��P;��W,?:�Q'��cө(W�$�\��]��d��D��S]n��r�m(NZ��2Vj5!�_#w��_}U����z�Ar�1h C.��h��lm� O��Y�K�dz�$)o�`�C=�K�`�W�?W��퇹/��r>B�������s�5!�L�PM�$�a��n����[��T G"ϱ����ծ��Y�Eq}BnTu�4�#��v�0d��K���;
[�W���=�p��c�ԙ��˰9J{s�����R��x��F6�&Ve}u&��I��BB���t@/>�Yߓ�����w�Yi�T�;	}���^$h���λ�c�i����C�1�;���Y|�`-4��������,&��8�~,��{;�Vs7�,@�A뀡}y��@%-Ӗ�=�Y%�nb��I90u>�$���I�����?ν:�l�Z�L1�t����ck��gGL���v+X�;s�Ysk��Gf;��*%�rF�$(�{���Ɠ�2�co�TfyK��D�@3��u	���m� ��UV�M/�7~r�Pu�)\�qb{����K!L�#~k��e��lk�R��o^���IW5���	��S*r$�e]���H��p!���f�!Z.�h	6%��)!���"*�,�tƙ�.�]�9���(I�{��zwhg ����+�ͯ�e⎌Ń����(y� �R����Rm#��EZ|�Ļ�h�+���r @m�L�YF%p�*��)��wd1?��D�lS{[�X>2���\oV��"�dY�v5���x�2���aQ.ȝ4�@����f��yP�wV���V�j^�)��6�ta�L�4Q�]j����V#�rz#�a`��o�7)�����o�{qF����R����O8;6p�WɆݰ��E%��>Ძ8���Y�73��[H��)�31�'�^����Ɏ�>w�o���}��ߌ�-G��X�I���ή�^��(c"ႏ�,V�g���6�EϷ�9� ��Yv����_G���f�!��[��C��֯��;>	���γ N��N�&�wEc�s0��}$�����E���A�ݞ?F_���z3�4�Յ"kd5;�`��)r!��Cc�\x �H�:DɃ��������P�Ü�+�_�CU��U�u����-��D�th�e��_� C�(zU�[N�
���6�?�q�]t�!Du~d{m_����b%�;�ξ�l��}��iu����y��S��m�;�*c/JD�%!R�Q��Q�ox�N�K��D$T�:�O0��B�$�TJ�٫�$R�����mK���s���j�0w�;�E�QL��5��QwK��̀ک8�܇� ��*��pc�����n��2�_힜�f�Qx��U���n��/&�Ȉ��:��r�#� 4�kh��n�%��Z(�[�G�y{Z�ECr�hڼ���Ռ��S�@��h``�O��-olG���^��1��`f��_�E8."o���tw�뮑A�}���^��-<�|�H��U�P����gv����Ue��)�9	m�)�@E@0P��s�&t�4�����PT�{y]��s��W�8,Meu:�ˬ	�7/�6�=2����T9Ae�~}�ZU�����wP��ǅA��D�ﮥ��:�1l!����
q�$
~	���{P��,\-��N�<f_.���M0�柊�l��Fִ�PmՋ�W�?Rc�����M\M]���A����i��K`��1N��8m�%,7��*��(_�!�]���Qw�1�<՜���ia?��M"�Ċ�Y_�o���w���޾��\���-��}M�SA�	=��j�Yw�����f��!$yW���d;�.w�E��gR�"�)/p���CQL�@��o�fn�7j>�l1��@OoS���˕��}f���9��o��P�h\��:�f��5��é4�DA/M9�dS�����U�
���N�Z�k]Bj�G�aݧi}���K�0N{�kF�.����QQ!���yzr��#ض�m2i��L��[�u�p4e�ɄټC(��*�[��(�jZ|�8�2��x��SY�q����݅qM�SqH!����[��Ҩ�N�w��3��/�~1���>���~�޾F�Vg�E���΁�K}���
�v�)�Wl�T�TΎ�?��v EF��O�Y:(w�B���yZ��I\��( �)K�q#x���zW�7c�.�Ͱ��6'"�n��u�g�`�8�kF7(������W�������(��wAߔ�Í��D�����KP�ok_Yk~X�:��i�ؖcƵ=m��aw�7e�lzS�����g�T$�Q�O'N��2�^)�����*����S�|�AMK�˙�{��C��L#%W:z�J�J����\��t��R�t��l��49��
����B��h+pQ�!��y�,\%NbxP9i�e!��r^1Yc�J�E3���CQ�y���f5Ј����Q�y��(·Ad�W;���X`w�N	U��-�¶�Z�����f!e��s���5�:b��(�v{3q+�C��Ouw��iP���m.�+�_E>��'��G�C����.ر�&���}�!h*���1#^x�`$ʩ�4K�����~$�Ȩm=�qɾg�����`Y�@��lS�-�[U�����oр���N:�f㒗�>݂�S������G��z7^Z1��n��Pq�vb	rN���.v�i�L�$��pDY���z��)pe�'�Xs��-^0#��[�Š�Q���3��k�~@k�������{N��Z���~��qU�]��E�,�
о7̨��{C�IN^-@\}����H.����Tؖ��&���*�����H�gĜ�,�����h�t;��_��\�3/��w����O�ʏ�皩�ŉ<��yK�m� R�����K,;�ZZ�%i`��<b�7������<��њ��F�S~6�'0����Q@�RS	.��t`���BݣM�����܅�����S�th�R^���t|`-l���[�׼��,g�7����xI���3;��T�	=E��+�w��$��Tn�c^���qN�>�\ ���ѐ�{j�q]/K�� f�zȕ~ߟ8��|�C�$��&�ۆ�h�?;c��>XJ�upK2U��o�ܖ`�i*�1����EQ��T�N�R_L�	ܔF�
~}�W^DQ�&݆���[��h�X{����.��![y�6 ���Y�RJ��w���1�j?ks�҃���R���NNl ��y&��o�z�w��}R[�ƻ��C>���vm���Vw�%y�\���J� [Y��P}����@r��x_>nFn��lAR1�Q��Gj>�U�p��A�=HN=�T���� ؜g��\75,Ҁ�@^G�B@ʘH��"��附��4�]s��4F_�Dџ���(�9.�s�
f�e������� �$ԣ�՛�X�摷,k���c��pW����}C+usS���s>X��A2�(4�>��Ж�4@*�C��=��v~h+��ƞ�\�)�������t ����f75��6;)��HN����>�MH��e�����������:ES}˻���?I�[Gi�'�R� �᯾|%��!���a����5�N���H3I3�Qbǈ\�r�Gƃ��/B��Ú��=�:2M�&_p�<>D5��'�8P�h�!�2������a������?
!W]8�G#�6DIC��>�l�C�;`��Rً;lᕔ���#L�����hjA��0%��F��5��U���I�(�3@4�Q��=5�.�Q��J����H�؃L1a�Zl���wcY ���UX,�@��@�Ȣn��cB,\���,���~��'�SN�z�)���OS�7YXse�Ǝ9]�b֤>�x�Jŕʢl����p��qg>�+����e�R�;4�坖t��S�k�5ˣZ�N10���6�� ��R��3���$�0�X��G�����{�g�Q���;�=�A�q��.��$E����Y|��T��{��Hq{%2�bc(���S$�7t|'F�y�xG8'L�;��DQ�,'��cl��y��:j�>l�je�������ԯ��λJ했W�����FZ�'^��+�;v�鹆Z&�|�B��b�IvD�0���xS?:V�Ĵ�D"uD9�~�%�ȯ��TFe��0jn�ܻq"�B�Q�E��D���G����g(H�H�������㡦roUн�u�Y��cU:V��{�Fk�V���̿���';ǖ�	�N���c�y3P�o�ˏ�J�n���y�-�{_X��l��g� �_�J}��Cj��]_����X=x���QK�f�5���$�;uI��e
o�<����\l�1�Za+��Ͳ\��..5"��j@��p��*�";�O���=֋Ȝ?��<J����� �75]#	LN^��`�[�ٿ�����Gh�����UKe�0n���?�еcS#N�����oŃFM��X�<x������>��h�fJ��~9:ı+������g�o����ː��O� �JczS��Eu2���T�D���<�����*f���� �LGN��$��{���K@RY��#�A]$�[��j7e�ϐY���{Ȩ<{<��S�u�褳�׾o����*�W��Щ"*�C��Ã�"Z�i�pq�&�:�9LY��?�Z$��{-dT���&���c��"�SC���W�"W�*� ��x@�a�����_���N������i챇#�������O�C�\V�{H����t�*KO^^I��>i(v���T�v��=i�^�r��5������͓��P[U��u3��5X�%�dnW��2���Ҟ�� (�m�ߖ	��>  %�9���)�6���2'5�(�*a$����W�g8�l�݁��]a�Xۜ�j
m�0V¬��򡷑q�+�����z�~�ʏ�9$��%�/���ium̞�G3�B%uU�����i�8BP�$ (����&8�WV@�
L��Ħ?S�M_�8�u^N;5��x���ue�R��"�&�J�l�{O�Z�2�/ԫ�a*�9�o�G��F��(�W�����p�iO��HO�!:�l^���%02�`�M	8���u��)2����WJ�m9yK�D^�qS����+wX9}��>��
q��ra�	h~ś�em@��W�LA>烚m�V�4����<�k�N����:8�Qtǐ��b���Xs�x�x�@���ںv�T������T�RS�F���X�n�_&�[��;𿎻	X��\n�Fk̪���ـ`����U��$�vgN'��A}�,���޷i�
U[�U|ͼ�7^�����&�e�)S���/@���Wq��O�<��b�8�de36��h�KF���lh=l�:��'$C/1Q�P�?�i�P2��o�#iaz���YpcLO`:Ij�� {c���bv9���@z��y3���h[0���ҫ|f�]�w��p5w��:���+�h/+���tfE�I�v�w����Ջ��}�}���)8����5��L��%�k2���ly���9b���N�[}��(�A��ؼ~�����i�r��l�2��ԗ���'먻G�a7v�ȓ)4hO~��΅�ݱ5d��ie��z[ň�'^��}�5I�4������������;q�c��JW����(�jr��:E�c�fw\�!=�X%��2ytߣ��v�Ȥ7+���)M���|��5Ļ Fq�}u7D���q��P�/(�N3�7O�l�l�h����a�7���;J� ��^�NCl���w���$�|��"��/!�k	2�������D���,�EN���	(F�&+Y�f�'�#97q���d�fP�����Zc̈́N"�醿pC����Q��G��K���S��[y������/�|^���J;2�=�y}r���V�Ǿ4��޴Qt�
k
��������#�5�!ڃ⸼��4M%��W,��/�����
OE���;�$i�E��0I�r*CՓg���gK��)��_[V5wxO��������_�i�����|TL����Y�<c�?�xz��0���ӎp4�5�.
��L��=)���>'զ����*���l��n���bN�ы����˱pt�%amUg-� 7�0�S�)�E0�)����L�J(��}�Z�����N��|ܿ�r�I�2ޣ\����SpAa�_+�m+4�x�&}���j���{YМ FͲ�Ov�U9�bʯ�#�rԻKv��3k�Ä�d��9HU��p�an܄&Ld�(% ��;qKS�0�y��&����^W�� �vC���(5��Hv8���ٵ�'�r���lPߛ=,�,�� ��"@_,�=Z���*�D���\�}J��J�w;�G��
܊��9&������(�����c���jxJ�L���m�����Msۺ$�K�%@5�p�F��ll/�]&� 4�g�B�u�՚$��TP�X�u�
	1�Gc�h�H�;*y�&�������i`m�^�ܣqq����BH�G�.�@�ۯ���[�mXYU�ɰ��w�(���I��AL�f�����gxOӦ��8i��v/_
3۷���]�v`�#YA�	�np���b���; Pv2�/��FΞ3s��D3�wD{����m�"��S�m��	��.E��q=�/��+��L��������'p][EE
D���P�v��\�����5Ui�y�x�c�mA�e�װ��k<c%	_�����F��6��t�(.�k:���e@dwE790�g;:�}
����2<B�M4�$�K�)8�:��$�55U6<^a6�Db`��l�%K1�j������~�\�]��A`˫tZ$��_�e��麴{�*'��Y�|<+��	4���RA���C�!�Mw�!+i�V�_7o���RVp>@��E��C���P��6���6�b.��)�I2@�%q9��+Hv	Q~�ď��[z|�����}�0�?�Ot �g�|�.T����%��Ti�"�)lT�<@����)~P���O.^K/�ZV��a����~G}�$S���ԝ�g�1��"C��M��(��t�E������L�����aYFk	q:$L�X��0ά8R��DX�U_>�(&��9�=;��P=��up՞�C{Ƌ�n5�K��Ѳ���@�����e��M�h�u`�h0ϵ��dp^Lz@����L���);���?�z]����LO��rK�̻YoM��=�!�f�_��b��2<��P�!s	��O#��A�����xK`H��>��]Wɍl&3�fS�e��O��&\)�^�-8�ZD��������!�iˎj.�)�w�z�
��C�t�'��>���H�\M��Fm��+x==�tF>�/���q�o�m��NK�Nꓪ�9E^/Ks����c3IB��� �~� UjƚM��H��#������:�����p���M�ڧ\����L�I�H"rY5��������
����1��Y��c��iO�k�XfOG1V�V��H�0{�s�g�_|^F��C�R� �u'	*wr]���rB�1+�EǙ�}�7moX!\c@H]M�d���`.����.�d�����ﴫx���	H�Fc�&�em�XlxVHYEB       e      20]��y?Y��76
4T���}��E���*R�9