XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���0>�Jf�3���^�S�w}@P������|>���R�˕47��@�&����	��:k}祖�ǚ <��. �(D�:h'fj�q�@�������ӏ������8�ϟ�gވ�����|�Q^�g���M���s2�/�֋W&$���Vt!�҉�@%�m|�RmV���#y�S��J&��,rD�/����Z����[�����闳_�yp�{1�Ȇ�wO�����S	;Qd=���]=
�(��8(~sS�����U���/vL���$ġN�$�J�nåt�~$��+zk���[�#�/�@�l}�{�͙���;}���${�m�����3q[�t�7���� �ϐ��s�yi����%V�u릛����g��y�w��P�^�*��,a�$��WG�5�;�$\��tI�'�����ƿs8JgsQ.��[���q��$6ұ�]P1�A��x��A��_�F�q����Xڭ;�LE�юy+Ҭ�wb�({dS�O�hzC�=��tP�:�-�>o�٩�i�����B�&g�"&Ra����������A���ל��� �/�j�rOg&���q�F�.�U;q��$@}�-�!c���{��qR�@�+�����|���v��҆Wk�NE�g��S)��K��#��+..Vj0f[�ԺE���Q�w�{˛�&���X���]�k�U�ڃ���)^�^۟\��"8�;���Bʋz`�_ͷ�����<�T���$��ܣ�O���<�B�6�iQ��@vzKXlxVHYEB    3b09     f80�b�ւn���a�|�7ɺ�%�_<ү�[�5b��y
���ZP�i�6�g ���Q^{2x�ߨܧΟ}:�f�+Hǟ��DA��[`�z�:�[������qLg8��PEc�㧀�'�ļ���_��ϊ�A����@�2S����� 5�Y����C��5g����RL��2ˎ�q�\h��B�����5�ez6�4[�ᰜ��)�	%[6_&!NKN:��8	$�V��?�1�\yQT����m�̝�!�̢��b��~�� l���E��r92uN����<Ie�kQ�9��*�,8�@����aM��ڐ�L,,V���9�/�7ņ��J��c ˂�~j��Z4�(�c�O>}&�^����|� ĕ_�qƝ0��~,�F��]��Nv,o�>�v��1aLo1k'��F��~Ap�a�����R`t��a�C���5�턆wU{ʉ�?�3�\��V"l�)���$U��\>Ӫ�8�zؚ͏\���$:�S�Ėf~�T�����F�r�)��Y#�'7�����6���F([%�:���<�:?��!ʩ�Ï�G2������T�a��n���Z�&�p�hj=͏H�?��Z1t�_����d���]q��-H���Pz�_~\�u�Fr��ߺF�m2v9w5�~� 2t�A�Ը��z�q~�1��2g�K��s/0�z�b?S���F�f�̅�S�ƸG��U��W���I�ś��^)(5�Z�M֦�=}�P��B�q�U(CI�ŶnV����$����4�,�͟Є����]�o�Yy�F���S�
?��_@���i�k��B�~U&j�+�tT9@",;�R�{m��#�Q��v�����
3,S-�J&Z)�$q�LZ�z�_���0���W0��y����4c�-=�1�v0�������oe����G�ԞkC}��e�lk2%���SgPP�߁!�݄&�,V����Vr�v�h\c�,��L��*<�œn�*���g`j�IS>a�)�\:6�#�3�b>��&q�˳Iy}mG ���P�<Z�K)o�	onZ.����lg0NϩQ��|��=�uvN��_�B'�������=.�fq�uH}{}ԟ9���������
��̽.��W!�u��ڭ| ߣ���["=A�PCoB����4�t�?�4�����܁W{H����i�bެio�׽@Bu� �?��"_M1�l�S��߳�v�7]�{�k�ψ�9<��JC����<���0�?�p��2�Rx�`�q3<RN^L�����>&ǚA����кІ%�ҷ��_�B�������<}D��)���e��p�i`q�O(�w�Zb��W�!��r,o0ܔ �0ؾq��H�L�M@�7^�b�^�݋ކ������9
3�z���y>�/�w��r��b�U��&c]THi�a1r{g�w�^D���1�I�I��c���U��8�GY+��� ��%4�T3���ډ,u��M�����PRM�+
�N�N��s�<�/��$� ��֘�	B�s��`Jz�T_��J�.Pi<,b.��8��傪"��|�ui�tV�>.��)�(�Q��� �ԐE����ܺ�M�sM�{1ϥ��msj�q*4�l�������f'������~vC&���ԃ�D�3$��]u=���inm�Fر�^Ϥ���c����Dk-�aB���uн%j���iX���SrMS�M[����a���n�ڠ���X�@h.�˿b���l�h#�D�'�������0��5)y�N�M�!�Ծ�m}�M�$0��{=U�j2@�+��۠�v��������xcǩ�z:K��dQ��A0�?�D�����(6 vO6(����ʌ���*��r�b��߶�Z���o�Y� w"�h:�e�+ᣩmEAF�E�b����~��%��[��/&e����CU���_TO�Xvi��U�P�bpa���W��"�>8 `�w�eMs��X.ڸ�D�X�v��aY�žbK��쎋L��4VP[�uX�H��x�+���Lӳr��>=��p�j���<Hl��JȺ���B�o}!�~X��>
�]s@;���\Mj dN���Qx{�~���іon���e�2�w����29��4��>��l�� �AX~�Y�*�b<��,�}@��e�o�CXg��!푢5H]���E�m,nc���b�PC�ވ���� c�*^��Wu;n�02Qt��F'�#��T��y�m�o'v/�
VD�z��o8N0e��$[��|%##}*�j�A˟�n�~	h9�D�]"9Hѡ�g`��J#'ɲ����:`��B����	ݹC������+�"y��S	��Z���3�,*�a�ѡ�n�c�'���wty�ƭ�la���M4ɰ&�90��z�C��!�Y�bSX!���V�N�6'[��)ˡV�^����n���$����$6蓢�^���ŕ���W��_p����x���X��zJ4���ه�M�����:֨�tA�4�1A��x?	�Y �[cʙ�OhY�_���M�,+o�BH��C����A�`�2�V}�?]�`�!&� C�/W(}	t�z���Tq�ls�Ђ|��^$��x'A�U$n��u��V��t�ⅼ !Y��WH����|)��EV��q�KG�P!���ᡲ<��d���e��o����������[�����0�����ɖ����07Ѓ'@;O!�TIA���R"u��S7�H�j�"������v�%"�Ẁ�P`Ql�;Rd��4�⁺�A��s�:��-��,n�M6��V���ɜn�!������*F6�t8ֵ?���8��g�k��o���=�8�<��m���ǻ����&7�-��QL~$E����7�p��$�Z����nX�!y�y�H���m��t� �8Ud�tNH��dk7'�2xlg14SGY��g��A��w`�D����s�%�	S��,S����~��?02�lBR,�W��?�Ğ,�	�1�U�8��BG|����ʦzU͝z[���a�����^}~�5u�u��ĒM`<v[�.�������j�3\�'�C�Vm����An�s�����omU0��; U�o}��8D�'D��<��J���Q������R@�#3���<��k� �v'9<u��~b<�W��N�>�9�X��ک��Q�;��XFBVn�=k�x] l��Du`Y�&+�ə���s�9�!B��~%�iR�Ϯ������=��b��3��s�%Y�"#G�v؄*	a~��	 ����u�uX�Op%��8������T�Gc�Ӌ��W~Ő���0-�G�W�I݀����\��R+��R��^V`㍫x��c�R�n+1��z4m� ��f��f����>�L��j>V��'M���%�8�S�z�-3��m�ay㴔OY�v�/x�y�W8�*�~*m�"]�HvOd�l#��.$�s��+`����t����|/������k��H?%Q��"��6�i"�K]fЄ��aC2���.ގ;�ۈ��l3g	�/�ĕ���ZG���W�B���x�V��j;5B�{�B�+�7����i����L����/$��ɭ�B�Z����@6�'lIG	�\]�R�f���/�ꔝ���Bꌠ���=������_�|g�z3�n�X.�-���e,c��1j���-����k��k������^���~��?��N.94[Rh�.�qy���GdO���I~le�{jp�ŻXi���ϖ�LRf�0��0�Lv��D�Ex�-����%�"M�+��.N�˽�[�9F��-�<�^6�ʬ��v�0�7<:����92}@Nc���� �!���C:h�+����� �<I�s��˘�2��`�KB�[G���t�HXq��qN��&̘"x]����4�}h