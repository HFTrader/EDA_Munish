XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bO��67�R�=}I@s'�mr
ن�.@�k�-����5�e* qI$=)IH1��R�u��o���0��/4��+�a�_��=����6�'����S�fF�S���Bލ����~�R�c��~D��}���� �Q�p}�cG˚�c�	�C ��&n)S=���ƉK�NC�ڿ]U^���7����:��%�O�0��D9Ua�^IkĖ��)�ݭ�Y��H�Ծ�N(��^��G ���q�E�i4�\}�Ek�@0��g��;E/4;��Q EyU�t:&܁(�oh��!X�^9��J�M=U�>�0A��uG��"��o8:��H��.7]�K.���l�Pv�,sz�C��3� ��)t�U��(h�yls�rß"EVƀf�c^qw�gK�%��ll���;��v:�_ЗnU���wƯ*���Ҥ�"�V�� $�6�=�v�����l$ �I�&~gG]V�H5E�Y5x�N���#՟���O�Ố.DS��5�X�j0g,�@(fbYZK��hA*l��f�?���A����ss���)"w�b͠��h�"��d��GI�OCJI�hU��L�x$��-J��3�ȄY�y����¢1?5 ~��{�<����(',ğ1֊�O�hUAp�	$��g����I��΃��W[� '#�����_�^f�@фڟq�쀾`�?�k���3���O�}(
�h]����a���|�_�R����\�U��N�Z��!�2�u�Յ�ǀd�ܨ�tK2�l8�t���j=��XlxVHYEB    76a7    17c0R�U�4�R�� ��Z*Ml�)K?�~r;�5d �ۡ����g��2���K�㸩�hC�L�O Aw�i�7��0P����Z��T,�@)�.�ah���2��^��2b<A�(�:��-��q��8h��`��O�g6��)�ݮͻ�ע 4W��05�~��	�z��v ��@}bZ"�U��+�o0Ϭl۹N��@D��Zb��<	�h�hv�?E�� �z	��A3���g�=���u`s�SNP"�?���'ټ��&�YYJ�~;,5�Bzڰ�DI
�3������hԏp~$�E��˭���L��]0HZ�/x܈�M�1�Hy�U������_���	��<��œ8	�h?� Y�hv��7��M	�d%��k?Α�7�K�+��k'[��+n��J��n�ha�vcժo�����F4P>��?A��.��~����
�Fx�&�)I������r��&�D��p�L�B���ۮd΋����0��hAE�--^��"�o������$��s��˕hC��i�������ţ�Me�t�sԌ|���1�`B;��G+tή|�ߓ�"Y������o[�(��[G;������k��rq/#�)��t���ѹ��m9[���}߿��L���`�Wᬒ�ق4eà`��Q��h�*�F�#��1�]��{tL+?�ҽ3뱪�=!�X�|��<��/��6^&����!�˪�Z���n �����
�*���p14�p���^�z� Hb��d�@`h�y��ij���A>��J�P��"m������P�}b6:q�	X�(r�W�ø�"�FY�9꧀��ÒR�2.�&��'��'����=
FM������l�o0�ؤ�0w%�$�sU���2�Q������L����I�z<.�eY4���)Δ@��h�䶨��~c�)Gd:��K�q�ŉ��!�j��8���J^�}X�B�(]�� ��Au�z�P ����\�K���;��.���<���h�����*�^��Cܺa�&k��E��g�U��Ē3ܠ��]KN�ۗP�*�Y0�H8�ݴ1�З�>���}���O���k��oO�4��+T2P0���c������nv�dD�ޙ_.�����fP�DԠ'V���WlSh�.+���FsB��\l,/�	-��\J��VԙH���������j����l:�����0H��zA��p�/ݲ�[�RaɃ�.�9!T��B_ʷg��0�:#�~�YA=���bqR�Yw�;$AN�Ga*�q�h�/�W���%\���D��{�̈́EQ+҆��C)���}��J� ��@�ɾ�jvք��F�ɀ�p���O���{b��zO���Z>�ј��yѳ
-������� 0:���񊞧�|�t�vsP�'�_�Me�nBdO)z^�7��]]{�3�و��&�;ʔ�Q�zx�����/d�t����R�_,�'?�(���9kfp
7��q}Cj��A�m�t���k��$S�fsl�H�6�����c�,�������x���@m��m�-A�<�ܞ�o`�~A+���I����<��4��ۣs�0��\�@E��'$�`y��g�FC�G(f|���aV�� Ц�7��ܨ V	�f	iI>O��F��Vr�J��RJ��~��*{+�=���b,:�54q��+Z�Dm�ޢ��@���t�$��s��^���)�yp�$�j� q(
���ɼ��~	=ZY%v�Ï��J��d���0���'�����s��ui�&x��;�j*���G���l3��"ȕ�������ҩو..|02<�A�%2�hYB'�Zwc� TZKS Um1����������˟��G���z�'��fʳ�Gp+�	~o��l~��.d���@����a�xhpA�] +�Y�a%�M ~�U+m�>Cwu{�AB�;�PdR�s'm2E�N�$;����7g3$�Ӣ�4�ĳG���n�y��?/������v�Ҷ���O�N؄
�qDkw�G�S��+ܑ�����D���j��?^�9�q�G�p��a0a�BI!��)��$:��A�2BYe	\X?�k0t�\%Q�򄌪 K
��Q���Zbwt��,Gg򎪂�%6Ej_U=Ӓj�DQ#y����d� �w���B�]���f�Ћ��o �8	;�f�u,=��O�7(%�Ĩ��������-<= �
�Y�����	V�>�ܿ���xؑ�[�o�50-T�ž�Q��ý�a��O���-�	X
X����*�i�)B~�/Y	!���3�U8�݇ 8�f��}� ���[��3f6� @�g�g�0]�ŽZKdm\��>�ݯ �'<$�'�1��u�d�3r��VL9
�gS��闦b���)/=�� �����x��5㟲���Sq�U�ö2a��<H;dÙ-��>x�պ7�+�B��%^A�,�q$&8�������_����4�Ӻ����jr�
��䡮Q��v�$_��vW9;㱩�RA/	9VaBY�+\���8X�;U"��_�X�!�6�!�0y|3k\��z
gQ�B����Jx�m���P�.2��~���5�ʂ�u2&��S�z9�c�9���y������4m�����֯5�X�t��o�'1��}�_��M�����Bͺg;^�~t�T<.lڥ�Kl��p$������P�6��EQU%i�0������braP�Ec,�f��60�Ĥ7��/_�dآ��[o�̥,���:�l,׷��hb-df�;�g	��'�����/U�	C\��?LGm�4��6d�
��}�B1i��Z�A`̚�t��[�-�t���s����1�U�fu[j�R�!l�Ii����@Py>�QW�;�3%A�Z����������-�{��7�R,�$�[Ka�����v�=^�5ńe!0V�]���tWt���o�?Ҋ�׭�씖$'�2�;��
��G���W��D?�5e-AڹI�P2+�x�(�}�G&;�ŉ�
>��ݖ����lc�Q��Zm���57�����9�;AH��y,q�c�`�_��,R_x��n�ϧdJ�J���:]�?��T�-X��'8�UNr��cS��ݰ��R#��GK�ܚ�	 +z��������H���G\� ��%P��\��j_��,�H�I{��]O,fZ��J�[�V�9\4��Hy��H�@�i>�I��JXg)z�nOo:�7l��]�����d�{i�_Y�S0�����U�����x������{�Q�w�L���I,��k�<���0&���.�@��)��]5�Y��8r�j��A��p{���
d8|�v:�HtS"��ԕ��\�H���Gz������z��V~%�0�?�e�(��F�7�0\�ù�V�nS�a�8�e�r�w~����^�����Ȫ�����txޟ��G�*��\v�]��$PO�U�L��|��^(�!�h|1�a3#i��b��o�̣ ��}�'�f�"#��������������?���u�y���(&΀^K���R��(�@LGW���k��h�>��r�QI����rn����Б��݀
:��p١K�'�i�L�0��\O�k�q��a���r��=}�s9���f����PW�Ė�Wo<.�g��K�~2�ش��mx8Q8�g	�t����ㅾ�G�!aϟ|&���i��eO���W�=�!Q#����� �o��ҩ��������� T,c ��O��Z����W��ua��h`yI��,��<�[��[�^��W��hz]�k�>(IO�����~?O�V��rˈ6�����s�}9���Y�E��vC8R����h�*�E��]�J���;�
p�O�Ů�����.�2�0���]�LA��_\�g��֌�Ͷm�I��#�������;��|��r^rHȌݾ��F�5� A=@@��v�#�2�B�"�2�I�|����gg�bԚ�Ó�e���PHºv�:d�zC��Z�ٻ���jE���3��3�p����(�18"�V]�'v���R���ylWI�$����g�}.���]��@^c{��t���_~7�nҐ|˥T���]�����o������X.�U�U�1����{b�2ց��^JE�b-���J�VX}1����'Cֺ�_o�5���8�k�����ęD�C��B���P𬢘n��Ι6
$�n�u����4Hq҈�3v��c��n��l�}@��d��9w}��a�����|l�ޟ�p9AhQ�G3���hR
�Joiˁ�K�4$%�.�T����./�ʖ �ͷ�Z�2�e�Y��8�|��Y��.Ւ«��TR���i5x��Z�~���A�?app_��9�jP�ˋ�k����Z����<�aV���g�(�Ш�s�;�q1�8�Iq�ۊ���E��n��f�8e��BC��Dn5"唑��sD��;����]���L��g�4*����6�<���o%���7�Ϻ(|ZO?����ǀ���f�]���%9��a0����$
�������m�A�3�|��*�)K�0w���H����h״t�i�A���ntD?UB;	��&s��"K0��)��'����	�����g���B�\ԡ���BG�G��n�$>�;�dl�% ���;�h�Cw!�R�vg���G���\Q�!d=3 �Oy�б�����Tk�hi��+p�h��4Y�T��jD�/�!Y#Tu�3���5�JS��J=���y���� |v��c�}��8�DpA\���JdM�����g,��5��볧��Hyz�
#���\FW�m����g�3�5 qSee���� �J�d�8��\�3EF^����XyIu�}�ޅrJ����>�����y�����u9�':�Z�w���'�;�Κ��F�nFIO��n�/x��]晛������/���5��
S�Uv�c���zV�^F��䇭����=���%PSCO�~�t�4��IL�@^�:]��׿T��h���'��h7�2�R��>�k�K�.�����>��'I0)~����^0U����Z,��@% F=MP���1��~�����k�bJt�ff��JTcf�!���TY��U�2�%�RM��}� ���C}�%.`����IO@j�f���k�F��"V.v\�谢��9��f��dK��W��l�3R��c	�yqnl*��D���~lby�OB<����Ng��^2Sʝ�kҪ�K,XcD?�'n�چ����K����>ְy�3-��p&$<jL���:�1���x|l�*���K��06Ʀ����W�84�� �.k%7�ȅ$��9��q�wV���p��l�6�"S��ta�����pbn�����I�4M�"L8tΝX�c��Q5�Ҧ�w����<�D��K��ik3#��0�����Ǖ>�Ms�w��Q�
�S	hLoL'9\PacZ+�P�ݔ�`�ݩ��)Έ��&��)P|G�}��@�_���z_q&R���8�����Ȫ��C�5�Q㩊���P��<���	[~iejK8�BT���.��J8 �*�5Z\.� 	6>'���5��̂�PWD��Mɉ�nY!L�ۇ&H�+eՋY��Gjze��uH�[����~�%i�`��죻2S!n�5H	��X�;m4���:�*�����w�=�U��XG�݇���AѐR��
�m+tS�$?f�Ro�������L������2�iBq�rS��cy^�1�V�P��h�b���3͗	�sFz(�<Q���o�p�6������P&\#_�{���C�]$t�ف�R�O{*s��Ʉ9���:D����n��C�m˻��ZFaw9
c��-cbr�My[�;p�u��b8�MJ�[���`m���F���g����?��22�͓4\�OY�R�e�cԊ��������� ��S���-P�N �o۩�/p�pZ