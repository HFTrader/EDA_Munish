XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ܣ��EZ(���ݭo�d��D|��ȓ�C�c�$�KH��R`0ݤ-"lr@����4��	P���T%}{�翓�
��p�ws�g@?���T�y����#��J�!K�TLT4��:�k"_{�A Z��pm'/���t�p��W<M��rCS-X��=1�`W�{G��hL-�޴������-P�Q,&�jilz���@I�Gy���2b�ڍ%r��#ś�V�:�I����|;�����o���I�|��}�2?���J2fÞI��2n����;]�7n�$w�@��T[_�gx�A��9��h�O�U�<}���4c��!2h��E�D�,�r��h#�a�*��o�V�V� ��v�\�U1d�7�1�,_aaȾ��!�"MKY)���A� /*�%��9��+ �`!�o�m���7a}�1ޜ
�"�JY��\��E%��mn��5��B���ۉg���/s�|;�d�k#^}�`��	�c&̐3���#]HZ�dS�1JD�T��^?�)�8:i���W�&ߘ�ku󿞅�4��ם�����w�RᣵnW1�D �׃�u�^Vh����oI'[}E�z���X'��@�'���@w<�^yg���In��>��*���)�-V~,�z/�n�"�9A(jo�ѥ�F���ܜϥ��(�eE~�z2@�2`�CQ<���9��W%h_%)�U�A���P�~�ɯT�H*wșT;���9ĳ'����&�sŽ#����Q�Z��Y���S��a[���XlxVHYEB    af5c    1ad0�C��|�^_u�t\�`EA�$�f��L
�_PV�zIད�wȩ��n�U !�9���/���DQ�I.T+�����K�g��o@_OF[�h�mX��[T�J��Nn��k�}��<l^|".p��zIqe��3�2��b��΃��T��!%غ�zz�[x^�,�+C�N�����IГ�$1u�ȍ庳Vm�Ͼh���x��z2x�=����M�c��~�g��I����>�p�G�������A3_ ]�$O�e��o��7j�w���Vel��-�@���$"r��,]p]O��"�F26pS���A�>�Na�q
7�cl���L��ן�9d�n�4��b[�2���`� E��%v?��`��)a/�>�l,�9E��E)� �#�I� ������z�-�V�͕y}�G���)]�D����`�����1+G��a�/U�tS���V����v����+�&�I��l&"2N�m��I�t1^���a��ܘF���̷��]���Tkp��"k#����?a+����"���iR$0�3ܼ���L��9��]����YEE�!IP�${�I����Y!�}��bl���7�fGE�/��8˂�f��������L~>�+i:��r]Yl�r��u�-澆�k�	yQ�T��[�ΐK�䳴s~[��J7�_!^��Z%�*���}����1�s>��SRB�/����=����m�s��&��ߗ��ж�2N6�*��N�Lc|\75w[��$aAȪ�fP�`����NJ��H��_5<a�es �� ��Kp�]�o�g�e�<�$����63�6�L	�;��k"�dP\����T8��1D�6+_��{l;h����X�,�P�o�-��g�����V7/$$l�ܧAR�����Z�i��*B/��S�����Hй�ֺŚC�4W�I>�ɺ�A�eӥy������&6�ۄa*a;��⊜'W9��9v�F;����`'�բ���
K��/��jЋG�u�����N���>�򪝒��]��Pɱ/��[��������.&nc��~ؓ��*�#�Mń!�l��|䅵Pe�< ׋��
flD�1��;�ŗOY�A���ȇ���L�\�!�g*j�L���\�Ld^�2�$iAL�B��h�����ɺW�	BoZ�8�2;��$��̳���?L �N�_�"����vDY�`;����C���n���I�2$���.�Q�bn�P�M���Mk�.��F�F�F.`g�Aԕ��i�B��<��������iG���6s��JKs�_�f/�Ȝn9Ru{����-p%훊u���A�$��LL<]��n�����b�Tk�|�34;qZ<Iqꅆ�JcR�Y�W�ʥ�b*����
g}�b�����g���<��@�����)e'�M]Sڥ@����p\j&C.��6�X�i�(͜v�$�FF,q'��Y���K��F[�:#G������j�5�����OV;T�n��M��"շn�=K0�oqz�1&#���B�k /c��2�EgP���Ց��en�[�eY�r�
��:�(�����Y����yݙ���'g��N~6�-��������(�.��a�3����F`/@���lE_1��`$�J�F�e�HApf��	�	]$Rہn&{���j��������"�6[-�%���+J�7s쫖p[�B�����~�&S���@ǘǿ�I8�F��&��Z)m��V7���Xx��e�c )�~�h��O�2�<��5��@2�4�U�|xL�v!`GK9�ϟԿ�����Ъ�ͤ�Tq�vLB'Ϻx��'Z*�n������;D&[��Td����$�X=��yB�@]�z���Pu�d3�O���}
���:u7{d��6ZG�v��PM�`p�|�sU�("S��>"V�������̿��8��q��P$��*��و��H�t^�h�>�:#N"' �9jspy�h'�`�}}��i)F��]�X���CV%g��3��G� ��e�
�Z���C��%+��6�>�R�Wo��xXw� ����و��<���z$�Z��2tբ�r�$�ӑ�v����=�@�~����)3����ĝ7���kY[NxC��Z�CS�7��R���0�P����b���5U#>��*��M���ۜ"f�'����%�c��?jlWLeV��"4��+�� ��Z(^�������I�,��F�%�1�|��>���p�IRD��G�Ӡh�+XC����������a��(�!,w+縵�>/-�d�Tmp}+�|�*g���.uc�;c��6�Rг���_O�5Q��kc����!k�F	��0�m�L�ͦY�� B����麸[( } B8u9T�`<Q�����n���y-�-� ������4�M�E�Ϯ��-��'P&�����e��t�Δk6D�(�y���JT�}"��pg>�&�S��� Z&��հޱB��ٖ�.�Z,�6s�ZO(�����r��HD-Ǎ�C��n�?JW�L�H��/�,��D��̯X:	�E������y���6�c}�¾fS��*���*�L�/n�����Η�_ݰ�Z^iiǉ:�1a���9v��"�ʄg�s�e��87������s���/�7�vF�I��ȳ"���h����`U��"Y%��M�a�ךgC��,��Q5�i�Fө�ņ=¾a�u���z�����'4ڐ�U�l��cG�im��V>�Ғo���/�-\D)�@NWi+0rg�]���d�}4l`��j*�l��Cd�0V��(��s�@C�)p,�+�u����
��b�&y[��AXGS_��) ���v�����m���L*�1}���{�f�V�Cj#*z˳ZS��ņ(�
k��v�;�r�zC�D���%c�<?�j��$G�lvd�9�pe�WX.�2�A-QZf #�c��V�Ġ|y�D?��Ki�~���h�1_y��e��C.j�Su7?j��b�Q+�T0`w�=��Y��2�t����}y��z�%T�	��ʧ+2�߳��|-�Y��EQk��鳰vF�xG��b��F��C8:\��\�֪�������W���y��%|�Uݰ?�ɋ��,�]Q�`�?%������I���W�d[�q�)9����{���k�^5&��'�w���v-����p�H�<]^z\����^�>���r��q��'�s�H�2�c�`�eό�w�"��/P_"��/I��'�4<�������^N�f���X0ΜB]}�.�G ��%=".Nƈ����U���* O/��Hs�˭G�a$�lKmn�é�Yi A9Q|yx����7��5$֓������F�8�����$�<AD3w-t��p��[�F�o���PK��-����<� SKT{q��y�^�p�뭝j���$0�Q�P��N�v�# ���Mk�Vo_��}��[��v�������6dR�����P/���5��+UJxqI�5�w���kI������޲H[?�$v)Wj;�e���#���G7?O�aS�V�����^�g����F������o���ͺ�&���4�r�R��K��ŏ��i]���w����M܇N�DߴT�QwzU���1#�^$��-�����J�F�~"p�zJ����Qulޯ�������_��7��Fg�Qe���^�6�q(��3����&~�?����e�t�p�D��u���>���	!���HN���{h�񒕝y���C�,��i��n� ��~�ؘ-u�+'�]5AH]'��˳��N���ώ��r�';�oH��۳,*�>b>3�Ҵ�?�'�W1K���� ��1�! ��>q�Q~��a���H)�G�f�S�߅�	��޷�x,@	6��8بH���Gd?����H���7��i[�� qFx3Kj��yWd�M0%�mڛ�GNt:���|�ju�oǗ�!)�r�d)zo��c�p-*w�)�"�$��TEݙ��D�d���)�2NZ�.ρ<��J�>���ԡu�W#��M�A��ߙY�.OR�Czc|dP>W+ߴ�:YqqU�W�@����Â~��k�G�����n׵��\�fa�7���GF��9��I���G�˗�uR���ڣm�8����*�2$��Y�֒���"��~�l�b�*3�����@��a>�R��}��ЊQS��n����7HM�6������}:�lc��\q<37v�y�r�(��O�Ӟ1�ko+�bU�5ٜ��i&��k��m��`�|����+l�E��C�U���O�N)���(*<����N�����uRWʃ�|�0� ^�I�����tԃ�Ƚ���&���₷/��1 �'F�}`�
^kNh��_�`���I*P�YL<;^��&�wAYކ�:C= �B߰��k�[�ͪ�I��-٫GU���4������عq3D��{:YG���Å�E��eԅ��j��9�>�Z]x�0��}EG�5���8+�ț��W.ҳ���Wl�w=�<�w��!T����������Ʒ�4oq�f���휼=�+g`� �����c'ʈ-I�L�������ҏ�ZGH�y�-N�G�kN���kV\����Y�g��h��:'{.?�#��9��c#υ��%TM{M�+�trmN���p�!V)$5�L݄����z��B=�(N�xw8��Fk��ٓf#XU�?.���(74S�w �zʶ�.lB������o��N�c����Y8$EQ bso?�����\����T4�`?s�Aj��Y��p��l�@-��'"�� p�Xѩ��!1�q.�Yc�<�T
��p�P0�W�o�a����[ ���Q�y*5k0c�&�^�X`=�ޏAf螘�W��|��u�!H�T-5�+������$f"�$�d@,H-���L/���L�uq��)AUƞ-�Я;�eva@J����]�tE��[���(�Q���u=�9p"a(
KOU-�8�O+P�����B�y�53��bs$T��X�_�Ky���[U�U�YM�H�ئ��}��v��C6��������;�e�Zǒ��}��y�a�'���Bu�/��R�D��G=��`�(Y~a"�Ȓ]:!ԥ���0����4s䜕�S��[b��04v#�y0�a��-�Y!����F����!�}��K|r;9��F�������7�6���f��� P�N�/�AE?����@�Ѽ�]��U ������>�K�Y��j�vu�!�E�����2l��eZ��X�f�n�S�6��Ya#�Yb�\�oO��R���"�ٳ�BedA��zԍ�:�g�z�"�.bJ@���/ŲH?ϭ�n�)����z�{B��6MF��p۷�0#	`���,�l�J���BM~C	���λ�l+���V���TQ��8���^0�;�r�����nf&C��X-T���ՄdH��NE�H׼*;�	�~K�jؙ�4�t(�Т<(�	������>٣,��B��.���P��=nq�bnsj�qF�� ���)BUC��e9���&|�Z .����%�t�5ɕ��I�/p��ԙm��2�@uqP��0�4&y�Ju�=�D3Q7�ʚ1��m�A��5D�v �u�xXbb�>S�Ck!x�`2��c�ڃ�&W�fUQ��~��� ڵ��@� 0�5`�B�%���p��bp�\�+�JR����\��c��~� �O�b���'y�	$�)��#�0��m�߫�t&���-�7����T�	\�B4*����T@���K'==^���ݙʎ�+1��l�șX�e��R?n��r)��ؚ;Qc�-��=X<o�CP!��Ҫƺ��fY`I�Ђ,�.?C"��J���%���T��Łʄ��0z�M�]��D2���:����\�lÍ���Ե;�ƮD�AN�XI?)75zx��|BfJ�5�
5�Zݛ�*.j@`�?6���1> iT�R���Ȗ�̀A9j`��i`��D�Y��21�
���3�mo"�`�%>m<�p/��֗�X�����	T5�t����BԐ���}6b��#+�-�&��Hm��@���c�Q�$X2����cb�v�!}Nn<y�%�ތc��,�;�G��7?]9[�s��~q��O_kf���	��_q�J�l�q���?g^@}��ON!޶�a����R� y'��R�s��F���������*զ���|l/9g��Z$����hwD���܅�}�J�r�#�g+?��x��8�FN�ط�G
ű�Y�g4���Ω�W���E\E=�}N�.��"��]"����.�'u{X��h�8��MG�^�����/^�Cs��4�X���9�~���vE�Oβ*F�&�)8�P��eAԒ/��8�P�N�����n�tZ��l�O��~9�=�Q_+R�|k��|�E �U��z.O�,w��Y��k"Yr����f�d2^�y����Ԩ��K4ٖ"����U�^0� FPF��{5`\�,P�`.��-$��[՗u�f'��l�@����`��($,�ق�f�@��!�7v7�:�Hk;|�
k�����-*��C�U4Z�o�V�UH����a��)��Y�a�V<G*I�fs�>�<v
sY1�O�Z������Hw�')��{{�I�j�,x�$}�Yf�(�H7�˓�h�Y׋L6���E�Wݚ;��9,�LrK�b7g�>�Q%<���x1uZ�*�����2_'Z\h�s2�NQ�������Yh$��(�v�h%Bs�e�R-�:_���;$�_�-���eΰn�p�����yx��n==� 
?��