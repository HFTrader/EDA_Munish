XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
\涡��m��Gz�N�_���#U�ĎQ`��U����\�LP	[��u�lz���������+�M�ivA�H>W��8-*<�{ f��T�PC�/��t�P*1��EE���ve�!5��E;��&�Q���i$D륻2�7 �d��>��Y����ր�A�� R�;�}^�<?(l*�^�<�[2�"k$���!�݅ERy�(̂���ʽ���/��ˈ8ww��W��'���L��}`��l� (�CQ���:	G�k��#d&�냩&���Ub��^� ��a^�=Au����N���er�A�O����������K/| ���g�v�*�1\�h�������4a��)��M�ԇ<��W姆�8�9�7���Mb���)�#�u�Y�*���d�ߍd()�-v_oMNBi���j�L���nolE����"��� P5���N�S�ԉ��?���J�����~������^`CZ���X~���$������V�ϒa��=?Un��
R��|�月ՌހB���0B]&>N�oYv��w[��|��u�BB��g�Ұ͌p�5M"{k��M6�Eז��Hw(�2�8�=G|2���>0/{��d�'�ɞ�KJ-u$m�|s��0�u �`�������?	m�~�&�ls&tB�bgk3�q�j'x,U�F'j9�չK�OG���)u���y$-E���������� 
���z�6���
�f��2�M᫯iRٚ]4x���j���y�D�G�"�XlxVHYEB    1ffe     9b0�r��W����1�ʺMZ�4 ���>��k��K�bh�B��b��
����	�<�b�Y;����o62�A�HL7G.z��#�j�������Td�����
�̪B`����MC�/:��]s��Ѐ��D4&���Bf��k��Rx![N�ҟ��ȗ+<���Rc��W�R�4�_:Ԁg�"w��������1��O �����,r��f��nQzȨ�n����� _g�pU�`-#qS,��g4~�}����;4��D��+8��s�4�Ǩ�dbOUl�aW<cd@|W��`YH��B5�q��I�!�Gxi(̉8^���.yv,�=B�C�]�`lw�ڳ�0C���!�@{4\,9�<�4�S#7�(�G���pW�Q���	wKW\ΈqP�����޸��^M�Zk;���D��L��������5�����0Ń��2�����f��2e�Rą���~[9)�P�ը�h��k���y�xGs���RN�4�_��@4T��{�ɍt+{��9A�p��4�t�� S}��τjo5-ȐQLH�c
R�O�9Âj���b����̓�8��0F�ɗ{�cɂ�o#����|�*���޽�ټ{�p�>�P��uv�_.�b�����7q�Ċ���2)H���\ㅙ7�b��/�.����o�	s�Qx*��RY0���g��z�/�����m�a�p΍���v��b�Qk��+��>Q��]ڥ�N�^���)�f_���52=��dB��tq��Qoe+���|a�C�m/�'�~�ȸyG�G��n��Ŕs���զ��T����H|�M����27�`�ۮs�.}�e��c>��}7V̠�p��7E��N�otU�*?;�q�%��,6�9遽>�6#_[:��@���5�[��,���^���oBHA}_�;l�N��r�I��g�u �?�#��Q��}���j L*􏪿��xP�pQB[���6���]�����-�H���F�Gp)�b�<&�2j��>�ZK�*
��iG�L�.f�AS=}�YM�z��M__a�6X�l�^¨����� 5��Y8��I ��F�Q����p�J�7���b/�\�;�F�a�X����4aR��!O'z[�s-]��8]��SoV�ݢmm�;=|��,�����
�	W���H��躺̰� �`=΢v_?Wx�Z�,�I����=x�p�v��c���A��'Njs TH`���E��'N�m�,�D��Q�}�%�P�P��]y��i�1̻�&��RY��H�"P�D~k�.B�Ra��:������!l�%����j�d��R�k�q��J���Ź����qV�59�#Os��C�z|&/ �\�V�U���Ӱ���Ϳ�Y|���t����.�T���h)��'�o���̚��X�,���sH� �0����%�)���k�M�bǪZ�)����rf�h|�����t8Ｓm���c�Qz�iQ�ʓ�嚬P�j)@�>����!��c�M�-��C8�%�'����h�9��ƚ�m�&"�fĩ����Kt�i���m`s���u�RR?ƛr/$����9�O4��c(%�_P/�z�����4��B��܂@"ͼ��DK��� <����������X����^M��l{gE2e��2��i,����� ơ�0L�8W5��� r�3�
'�S��J�@��1OBRFy�9�Zz�]'n�6��>V�����~eK���ֈ.����r���ѝ��[� @�������재~��!@�j�$ =��+��Wce�{4���(N�PM�X�!���v��EpX�fLF��1�T�`@� VX���ng8C�2�z㶉b�'J8/0��)Ukj#m�������L��k����������x��s+�Q[�����x�Q�6M:q���q� f�\�Hk
�ɑj/�.)��&�|E��:�Hs���Ma8����n�t�d��o�.��@�)�-���X��N���N���\���7��(�Qr�1=�	j�Ěw^۶V��݃f���������8�7�'&?�.��wf��jO,�T��w����FbO%�b�V�c���������؋l<���x�^Ƽ�? ��H�6/�knޫ���wB��} �y�}9�vZ�:)�0��pcΚ���镙G%������v���"����	,�]5QN�NO���K�ՙß`4Fޫ�&���i�l���%݋4�b�=������-��Hq��T�aڀh�f��m���ܛzIUyԙ�{Í*X���5�"/��*�1�j�Wt&�@���Y2�e��0sdd�c���"�9_�(Q����Go	#�Y5��WDH���HS"{��˧�7&,޽i�gj�(�Q�#76.N�'�XA�Q��>5K���`&
�]�0'/��t�Χw)2(6�]_D�����LQ!:MG.�c_�x�d��h][mv�ɐT��ȓr	Px4/Ӆw��j&3�"Κ��