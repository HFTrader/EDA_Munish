XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��wEyj��h�J�pױ�s��r�aG�p��k": �R�gã |hm�(�510 ���u�<�`�"�g�8����=0�S� Tsٍ�w/cr�+��n��<�3ď�w�,25(�Z�<x��e	Z66��2Vz� ۽����Yf�����0�@�}�g��|�I�$#h e���~�u�[[X'��-,x��%�^z7��2����4�`г���C]7I��	2F�Jx�b]�Kcw�e�u���\K���;�Yݟj�Q��M����|�H&��u}w�ڿ�L��'����,�����i�����q�Z��1ٖ{��{h|����-���?}���k���?H���v��G}�������Ԥ��S�c���B��	�N�#g�w�;;��O9����@�B��t:���'&$_����q�zB߹���9��#��tA�I����s�Vn�>�~�iF��+y��&,XAI����� �W��{��f9h�)�?���dT���%3��듻]���G�&�l�2�� ���פ�T*A��il~v����&�
z�u`k�1�����1m@�+�e�s���$��u��w�Lk��?J ��!��E@�?��ޚ��'Č�|�3�z��%�(���%��'�#j�&������V��2`�������ˬ���ؿ��g�Q�)�����H�J�O��"�ُ��,��4�9���lOn�0����1C~�\--�A�����q�G-�ѣsH����fT�@y��XlxVHYEB    3fdc    1160l�2+?Ā:�΍9�j-�i.^�)C�g|����w=^9�̦��!�ʬ����jfB��t.Kԏ')%����d=��������z'癝 �J"RRVV5��j�钥��\�zhu�,�PpԿ��H���u<|��p�_-�ţ�7s�M?+t'g<2H���X�xۋ$� cȔ�$�Wu������N�� /$��j|��o�%,"9��3��s�LD���s&�Ŝ�ϛy�{��P�v8��ʻv&ڝ)}�a�I'e0eQ�~��E������W��,̨t�S���{Ho��#�Ś�� H����B����!3%:~�w�'�Æc��=%�Qp�Hs��z�����?<Q��<F���n��ڀ�d�
]�=�sQ��	��C�t�xR�I�P-+k�B䛄A�l���*,������X�,N��;La�R�(|�^�uC���]�I[�����V�vʏU��k���[#�8����� -V�m�oƷ� ��#j�~�� �s�m)>բZ� I8��~�M�Ro�mg�*�uv�@g�@`<�V���$�J����eM��t��,�X���>Q���5 uՂ�b�zK��G�֛Py{��g1�7�T�C΄��̯�#�<`���0I>_�f)W��Li�/C1���o� ؗ;�o��%9&d�:�ٕ�!��D Y@ hS�O^�����+r���_b6y��� ,E�q����M��H�Q�i�\ ��S+��=:356A7����^	�N�48;>)8�S=*�/�Bj�>ۿ.tB�}�7ȿnxuI�F�)X��$�"<͝�Xz	t
W�MYw����;�2(�}p�h��sJj"/�,Q��ٸv�+���,H��"80&�IX����"�ݜm֘<G ����J�ڤ� "���h~�:���K��!��ݵ�E���R�B1R�S|���G�_�a�r/�ރ�6��F����e�z,*�����|�Ě���_��u��h�D�������:��ښ�O����k?��=ӫEU�]&�`�5�^���;�_=nwn�)�E�-E�9�a����,Ͳ6Ά]�2A��|�8`�w�V���@z������A$k��Ym��ys�L�K:0�
��fU���	��	��)��&.�"�MCY/���ܖ���éHh|������M�|e��]&�~�!��p�9b��f� ���^}h&M��Z,:�2-�%$�&C��De#�4�����T���f��_�@���t�yi	�B5��3�Y��61�Д�Q�h�5�m���t���a%8rVAC��B����x����T���t�S3�Z"՟,P��>���6�T2�#h�;!%j@�`L�FOgu�Ď{���esg�d�n�UInD�F\�I�8�/�{�C����9؞��U+��A��&��%�ӝ�uӻP �G�3� ��������RđRj�j�y)�]����3��Z�,���`a�A��:�ۭ*Du��2���5�,�=�=����U{��1Xu=:ųl-wR?���|k%�an=��7��%�_�\�ځ���ҕ����E��Hk0"��su��<��"5��]&����ߘ �4^��g3�:���Q a�j�U��[68���/m���7X����*F.��w�7�0��d� I�J9����]�T�&Ǎ;O�������{���Cx	��r"J&��=�s�_����g%�Q�&�B�Q\�R�����b�DI���Lv����B���Q2ؘ�J��"����X��5סs��~W�v�@�������C���o�����������b�����V	&��;��2���=�a4QM�MSZ���!G?*��� f�S'��O�� ��pU.�,{�d���dp@��*\��~�X�l��q�n7��sK�6YK�j>v)[� =�w��_=) ����������{��q�0��	� 
_���:�d̄0�V@����Hc7�)5���OE�h�1�JIz����
4�R��|��򣉤ٴcO�C�H:RCtƀR�<i�P�������_�0�du,ᴳ����;��ޠ���_���p�l��~/����`�*�Je�]pو���9�Ko�B�d�Ƶ�!���H�1k���2yB �]4V8��HC�~�ᵐ��U[��j����;����,eL��&"�r{7"�l1&ڛrHz|���z n�1ȓ�'��8%��������T�<y`�yV����U=-�"�:�L��9�x�Y-@���?�n�Ć�<}���Ԫ�mU�gt)$v�T�v)�Y���~8��w/�Ǳy��=	��9�f}\ʽ+�����ȥ�-�OR����X��i�����+ݏ���?Zӂ-FG�˖m.�]���)0��kc�ӧ?´?I�A��-X� Ou�/o,�*c�e,��l"Q�^0�����-�h
��ﾎK|.�-r4��͠2/��~�55�0�F��ō�X-����j�A��^O���S?Bd��"]UŔ�*������9�V��c��K �D+vkf�!�^|O��k%���� �w�����]a켐�D���������y�Sbwg,�8-ro�o���9�V8��jZ�:�ptg���#D@(���+)8?5�Ӽ�k����N���7�+�!
)؆7�R�Nj���*�&M�~��`��d��80�Ni.N�;l��Q%�<L�OX��g����u�_��K��o�b�
g\>P�+���Z@�\%)h�OB�O��~/�,?;����n�<�#[YJE-Ϩ�/9�9��%�y�����W��~j[��'��&���D�}���/Wx�:�+�] ��H�࢝��4���A�>��xm~ϳ��WC�ճ#H͋k�k�%�ޚi��C�X>!�e'���K]e$���u�X	���+ƍ��� O��f��CG'�SU}��4��7�c�ڄL&g�ד쩙e+}@�H}B\������b����|�u%�49��u��͗��M&��0����n'7�T&L�-��-A�	ƻsrO�����3��8�hX5L<id��ޏ��㷎EU߲7ɥ7��Ȗ���=��2�f#7���lb�r��h$�����1J�����T��e�<��
�0��>�/�1.��r�4)���_���!�W�r�m�|�X�Ҥ��u9l���ۭx&�>���(R�lʽ�o��;`{��(V/�f����A� J����>uI�3�&�iY�8�'�F�*�pMÂE�� p�䀐��e��%����wO�7�&@n��Q`�hN�y�p��HY�����"��qt�����p�
�ܭ�f�	l�n�N��F�A?�D�jz�W��H���줧��V�?I�?����t����%J��[:��^��v���^)��2�����F���=��B���$�'��(#�
A5�I�n��؁��O?�yK8���D�����A���o�oѮ�~�F����
Z́��yqB�=�{�XcFj�=�!f���7�?��:]#�\5���D�7'�X6��'��=��6Th����K���B"�7^<��/��:f��l�]�+<)�TJ�-��6����Vg[;��F��mpK���W]�erq$ȭ�Y�.�1K<�JR�Ή����^�`E�ǌ��M��e�B͔��'�rQ"H���Fi>��n�91c`�z��&o��ԉ�֢���j�B0>S���M�l�;��D?c�Wc�-f�cp�Y$W����y�K�SS���#nL��Ik��(A0O�Rw�7+'��JM|��`Jr����E�������}���P�L����E֝�5 +9E����,�`ـ"�n���Q=�5��]^jx�;d��	������M�K���o�d��w=�ZH,�%C�~0���Ulި	;�9��Q���S��&N"������ʒ��!�U��W����:�P?a���[�$q���0�n��6kٛp���+����I�.Ng�O�U:x�����<��|#�j֫�]W���Z+��X���b��	���H%��o�nԳ����"�_ߥrL'?��ҹI9Z`|�����J^�#�SE����C����ڠ�؃�{M�E�H�G�"d{��S�e٥������~F�,a����Ʋ�ms��H��$v7��Sc�G��k ��S�M�R�#�.>�K�l���Q0����it��3{�q%'�����}�i���^����-�@��j<A��m_��u#Vϱ�QY"o�Z��	�@������\<��V"w����B�y�=O��r��d�b6���Ho�D���*갵%]�ۅ���E'O�,�X�QJ��2��ȶ����3�"Td���^�nK�q+U��y.�@��~�'6&�W~�� ��9]\ʳP5��DgJb