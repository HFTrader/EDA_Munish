XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���8�X��Q�M|����ޕ�	���_V���%\
3e�f�{��F)[:�����޶7��^���^����.���R�:9�Lԑ�G[x)@��89�I
L����l� nh�s:���X�K��L��(Zz���z�]C̸��<:�Hަ�N�]�TH�]�ߵAku����s+�{�h��$�M��S	������E:2���f���.x�����Iױ��H�A�@�@�%�8+v^/�-㐸�g��t����'MY��nהA69�`Q:Y�����F�e!o�᷊�ȑ��D��:�`�?���ӘH�T	�s��tr��Y-(ē�-�-u�v�E8iN74<2d"�Z�l�@��&F�-۰?�����u�B�V��Щ����:-�R3W��,�﵂���	�{����k�)kwM>���6�`>�h��º��$FqQh�� Z(���ޑ��`��m��C̆.�0�RG��#���69�_����?=ws�lt`��A��v�NI�v�1I"�_���n���{:�wB7�x!F������l6��D�o��B��X��T�4eR3�[6����e�u����b��͒c���h�{u2(]�4K�[	�Y���f��D�z6�	t�S�] 8s�����x4ͱ�R'[�(�p��������r��]^����Tq~`k�Ps��h����s5���o��{w����qå�͆h�X2X�G9���J��'��DU9�)�>ڔZH�PNw�.�b�9 .�����߂��egvWf�v��ٚ�XlxVHYEB    29da     af0B	k1C��߁dE���@�J�`[���T)�e��eJ�D[P�p�&��푮J���I�ËAS����t@��GRV������M���
�iƦ���@�6I?���\��ѥ���e��)!6
b���[O������@�^Kװ�ߩ
͠�����o7k��{b������F��r�q�ݽ�W������Ԝ��m������v#5ƭa��Y���_�K��4J��a���+��/����v�~L
W�Z��=C58�Ky��X�l���l՗в�E�ѣp-��k��l;[Ü�"�&_��l)Mt�����lr=b/JE�Y���}��
a���h`�k��s���h.l�Z���m�Ƒ6٤��{�D����#����ɝp)�t1]�����/�^E䣄%�>.gvt�+Az�(4��c��3���<��{D=˺�����7
��q�^�^$>�:����e��sK��V�!�w�����{$G$���T |�?KB���<��9�^:Unz�7��~�7�J�C)����
�a"8�f�wW�Q\���.T
�q�a�"��>"�X�{縤ɟ�	d��I��(-��p���g���ś�ڲXTٍ��*��j�+�	G�SYq�8Q�=Qx;£%S"AF-�(��ǈ("�>���sr4B~7�OB|��
L���	G<Ms(��s䏊x�A��E���w�+ڑ�3�I;��B�UZ0��Bv�!��Ÿ�(N��aOJ�ڬ���}�����#L�ZrZN���~⪉K� �I�y����=n���._��tư��<}y� I��blQ��	H�Ph�̝W���S��wg�9Z��Q���}�ôWi`�0���:is� �UE��CX�'Hf4ӔE��k�uC� h��B��7�\;}���>�ۘ��Q�ϑ��(y�C��Y��(s�<�
�y� 8�@�?%�����c���^��5(��mD^
4<1wY订vt::/��S���x �3��֤����������A�����7Nz.��{ĳV�_�ͻ��{e�i���'20�B��,�8 X�\I2����&�2�K��쾯e�;�<�T�����7�%/z%��Ir{$������W��3b�܍����_��~��;�v0�u�V~��i8����z��}�E�[[�)��1�^�����|x���7�_�5CH��̛���֩t���y���eE��Z.H&?���3�]�3-&�j���hP��0:��7�#�����6m�,�41K��L�I�j�OeaoAM��t#z��r�m2Wd?t�Ҹ��-U! �+ʥ(<P�q|�o�(��.C�B����G������e����� ��`�(c�޷%)�k?#,�e�I�p�O�g*��|��`��h�ʟ���@����hm�zd�>�������d�۳��?���m�%g���.�슈��-�g�Ã��'��'�%,���5-���w���Tm&�r�@�i�o�9��v�L����+�٘^"m��p�&�g���Y4M̟V�,��P�&T,�@��fZ��%�)�>Q�XUӜ2��B���1P\��`���a�Є~��^�l���c*����3�=uB��#p)�
�
��]΍G�|E��i�}Ê1w�l|����mǠ�s5m�5���\tC�Ȍ�h4� �ܫ`!d�������T�
�+r�R�SDLu���b0
i���3XxI�u���V��~J|K��;���
�\�Y����+'�6G�t�a�M'J���o~��,_����R܏�:X@7�5;k��_�M�w�i@Xo��3J��P���04�Ԅ�L$�D(�gW`�Bc��\U��b�~|c�� 3i���y�&p�/\{R��gUXP5X�H'���aJ��i�ͬ��C߀GM	�����)Ѯ�w��E�E�_gA3HYi;n\�����ڐ��*X�Xs�F�ߝ1���5�ϫ��#��(�?�<�+> s}n�!�:o��s�����˒��?���o��N�I(�$��Ot-������r��W]�41�0A�ֺ�AD7��.<���d��\���n�����3��܃�].x�9t'�D��ȫ�20��f��(K��vߌ�퇴A����w�4smzB6?�N}lz׷H~�#Q�Y������|�ʐ�Ъ�x���&m�y��gm"aV����W(�'d00i�3[:YC�N�: �1b�
LD�
�dn�dGHpu��&y_�2��GH��%��p�Rd���	�C�������gT��!~�آ�T&{<z�I<]�����-J7��ۙ9�{a�SO�!׷���g�Z�8}Nv�g�}�#KTԶ����P�Mug���s�%7WS��d�r���v��ں�����3g8��F΄`YZG�9T
p�9o�V�H�.��۞�{\VM�x�٤��9ߣH7﯉��4�����rB@N�ił�.r�;�T�K�����1pR����$��d��Z7��cf�#f���ao��'�@�aH2���_"z��I�h����`ͦ�"�g�]��d��;	����MM
�B�	G�4B$?�+P����MW�q��#�Q����oM�l���g?��i����N4i"�����\����	�s�4^GG�h�䧞�B�rSD�k�F5��g�n��� wm���Z-�y0���Uw����t���+� ���}%���N�bN.T��`a�2@Ǘ
œ%��H���~�t����X�5b�n�I��n