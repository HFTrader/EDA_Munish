XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{����N��Ɛr(����C�0|��������
���]?��s�HF�s��ޣ�@�m�հ�� �,t��K;�.�����y#�kw�1t��"�6Yt�t�/	�Q�#0� �^�
�:�k��'VPx��9�J�}0�4+Y�fl��;�U�ݤ�]��ø�}j������Z�hAveHk���BH �,���wh P�-3�_��v�`(Y�zk�X��p-��K�}=��H�e�Ӥȃ�o��u�&���G6�ƃ��W<=�k1SN
g�H�7U�}��jN�d5p�<.�)�;�����'Ww������&�
��b�2Kә�i,|�	�f��$������h�xK>I�>��S7i�����A/BЦ�\$*UOP�����d�Dq��:Z�J�Œ�~1��!ٴ��W|�S�;�Q���6�~"9�zq��t�v�Ti8����`x'��#ާ�9[;�3ko�a�ha��
99M��$''�6م�T�.�Ė��"ē9f<K�If<�Q[��rי�������Y�[���7�$*�c����6�A���k㽵��:��B*��j��0#F,��|��øB�Oj�rj��(��nb�mA���jg.����:ٲX�#��Y�z�8��tnN88SP��Y5 ��a��5���O���I�Ȼߍ{́�k"��,Q�Q��qwM�+#���� \�3i=�]C���Z��K�_��K�c��,�K�Li�z$�p�U��!&�"�>� 3`4�j����k�XlxVHYEB    9732    14d0�<��NjXW{�	�Qt�R�8�ͧ<L�f��ẕO�Lq�>�p�p;e����4sLXh�'�kL�Yȳ��F������5�g8��@4Y	Fu�������{��g�� i�1݀A9*)�.�sǓn?$p6�F����)�N��a䝳w�u8/H�r
��i�g�AHy���V 8�|����L�sX���Dߌ�x�5o?�ؕ�qjPN�r��%ơ��F����;~�_3��3(��|��j"��GC����������u�f���G���-Q�^��N�фpP�E����Q|w���E"���A$���v'�>�i�
���;{z�e��Nn�w�(��Rȍ����c���	�ȫ$XL��U�A�H��w spic��Z*9���^~�� �_�3�����O���_w���&w�љ��*p��e!��5���:U���wI�y���@;<����^B	�0��,;y@7_�|p�����P��i<����`}��T¹eX�͏�S��P�7�r�7>�҇�ؘ�RekG��fЌ3}�L:a&3��y���]X�}1?��̅c�c�ݠ�\�v����)2�I�����q���m��؟U���LK_��q��0z{����Gڹ�����uBq�O�.�vRMQ�v��)�Q`���c��)E3Q�`��l�k��r/̤}Hqy;5��>pQ�̯)3F3���y�`�:�g!��x�"3>���G��HlXņ���ۛC;�f	ZL_,��9MH�n&}��O��u�
����'���(��B�_�e[xD��'�JW%ϣe�'�F���2ĵL�v4�?����l���;Hv��֊��(�ɷ�ϣ�_R������KS�nXځ���ۯ��^X��?-e\w�W�g�<:kiͽ�knM�n�ݥp�	d�'Z�:���C��y�c+c���&I���g�r�;��z��t���>�d�t��s�o	��2��\2C�L��F��$��
����P�?�~�9��l���6������p݃�ݚ���;Z+Z�qjC��g�R�&��N,H#��}�̟�V�~<T4Cj���B���s7�����y��Wz"�pz [����1���	�\sg�W��rVW�dP��ޖ�ˊ\\�r#Ut=����Aqoo��Լ��΅�h�F����k}f�	��a�'n�"u�G[��:G�ݷ����b#��6�I6b���al���*�iW��qf
4e�Kt;��yt�2�؄YzP��u�6���:�	W��V ���)An#_�L�nJ��`���u�����������3�[D{�Ӈ�G����f��(č���f�8Mw-���\��K�M�q����1�~���@G�����3������%<#V�a6��VhōUgy�f*ߜ��0|\ MA����U��(��Q�׃��ze�8q�uν6ن̍��.<�c�c+#5�.>%Q,g�F-�v+=q_�.��*tCN� ��lXbmgO�xV��r�:�#h�[��v&lf0��c�X'���b��ƒ�{�ۓ���ݟT�G�Z2�3�k!��R��oZݯ�9^֦��K򲜲ur0���������yk����c5c����ٟQ��/�5�������[\t/��n)BQ;��^��%$t�f���˓l`�(��z�~Ǔ�V��,�̦K/����O��X)�F=ť�����c��i��.6e)8v�\i�0�m��f�̔
���%k#�|t�\M�IԌRf��U�6�]n{�)rB�|��k��Hg��tWob:D�~�o0�3>P��R9�����A�c9��9��q�2��+���rQ�b��\�׸?D(�h|\��W'G	hP��;aB1��:T��VC�A:8���V �%qy���l��F�P%���,���*k����A�^K�MO��)�N����n	j��h��>�x^���2�\A���z��{��V3��j`�R2�J޼�:�i��h.�U*i�;"��E���4ȗ����)�teqH�)�|��&Q�dT���ɝcH}�c�zW7�*��� �5�֥�:�zg��(%��RG$ah��u-!��z�N�Y`��+�Hؼޘ4�T�3�c_��t"���p0o�Qq��uUf�J����҈?�ӉQ�(7m��w����з��ej��AuC�ė��ϝj7�.�<c�:�Y���Ц&���lf�ʙ���9��Tg��1����2)���&�� 'ڔ\6t��~£ ���L�Fe�v%Y����u��;s � ������n��9V�F��Z�=r29���Ñ�x_���q��wFV��Rf;L^oq�r��p_��pm�:8٧��ρ�p�QA�Oo8/4킷zT,�'qOj��2%NL/�)u�-�~�3�瑕�=Ī����?��XQ/�]UX�]�c����r�mm�n��B�>��T��c�.���o�e�f��%�9b���S�,�ފB ����آ����u�; ѕU�4���P}]�����'� F���5a_��+y6��O��]���s����ܳ>Ùyz�R��	�%��d��s3U�GNk'�I��ǎ�]�^�T�i�S��X|A�j�d������{����ڽ���*>�u��g5Ff�z,6.����;q�ghܻ��H�L���z��5�R3�* �e~�8"ǡ���=^}H/�MǪ�n9wxq��7��az�&C��U��c�|��U�E�� �ޥP��0h�&�{�N*�ٸ�C�`��ʛ/;�Ѵ� � 6g�j�8Dj%\������1�W�Y���޹�Eդ����|0��d��k�.�5�D�0�/�>�b�\�M:�W,LGT���H����{����d���K�j�E��

L��2���=s?�D��b���%�O-�p� � �(s��R AeC��B*Ԍ,�L5�݊i�ي����z=�]R~)?ۇ��I���/���&�c�G�H�c��B-j	y�B�A�3�s��[	<�����
�M�k��*��h��t��Wk$�$�5����	so�TO����<�P�� �`|n
�%���Q�=eA��-+H����3�hy��Go����a�5-1����q�v����ÎF�זD$/߁�(f8�| ґ��^I0��U���W��lSyė��*����(^��}�$�[O,��3.���xxv(�l��S�������|��#� a�:��T�WL�m�x�Y(��_�-`j`�`n��Z��#6y7�9�	��d���щ��	0lo-�L�CS���f�
T���-N~��ɤ�7��� ��ְk��1�6���W���&x�K>��O���T��'�����3� �o�jw���L�Q {N!rFz�ZF����b�:�_�p�o�~���!�����^&�$��K�"��{�GVϤ��߫&��!Y�;��v�e��W@m/��I��)�I��i�[!�P�>Pa*�	��j�GW��G��C�K-Ӊލ��M��p�'��F||@�Pm��-6�n�f#����߶�-y�y�иOX�8��e�C��|��y�3z{e���b.�?d�w�h�}��������5d��vU������.@$fI���K
�.�|>�3����i�#$ُ�n�8t��kW=؏R�k����[�h���᳔�U�T�7�v�u,����<�Z։���e����^��M���l=^�?��YL�
ા�cΚt�u
�ݾN�}**qҚ ʝ*-7C'�0��DF}�ta竘<�b���2[��{2r �|�؜r��rЋ�mcax���4:��eTt-�c��g���@� �j(?�l��ӭv�YԕK?����-�wxu���2wq>��'֗���q����d<1b��.��<QY,&ˆZ����v�mґ �)�W���'�dM[	%	�����n�ίz�g���K=I~Vn�ٕ��b��y��C�&&4W9���"
酭��B��̃�k<�����l�T�9��b�1�`���,�n$�A�9�{��g?�YW,Zr{ay�xJ��!��I�v���b�/���˷�:Ծf���@M���(�=5��3��Ze�?0��3����EW�)��ZK{m�n��-���EF��w��M�o���㣜��w�g� "#w��*{�FR `\�M�=��*������v�(�]!��3�+�c;<0L5�2j�� ���c�+ÈV1|�'�@(%��Z�衤����2S4��D��iV?����X�I����œ �<r����..��>	c��U^0�R}j�x)�`R{:`��D�y}%}`q�yC>ғAr�m���]29���̨v��YW[*����n���s=j7���(�+�r�A�eD:����
���-xA������|���:��B�ɭ�	��MZ�$�;#2�M��ᱽ��Geʏ7�pdIj��P�Nq֢���Q9��{��aDW-�gɭ�����"��4$�j��3�I��?��P	�1�8n\�\�\Sk^@(�kk?�'�y�ð�H?�iF�T�d#�����s8�'d��Q��N-
יʃ����NZ��J���%��JӾ��[���z%���OfM�� ��<�D���*z���ﭰ��*��%����($��I����>�O4��Y[~K��I@E��#�l\��ۀ�O&4��S�(������K��!�~��{��l�n�$Ŏ���^q>}s��	�9������Ba�M���H���7,G��W��T�����Q�V���w���[@���G��ME�4�g�_�Ġ�j������R�K��v���>r�e���2fW���k��<v����!����z�'�E*[B�'�~Ӎ���ZD��n�m�w*�t0�{ߎZwi�#]�!���*��[1���4f��7`���Կ�=H��LoXEb��w�������z��Lh|ϐ�@��B煟-�^M �Yg�}w�_��%1-��v��^8,�\��{P%ݯ8���i��
�z<���ސ�o�@��B0���`6斔���pΎ�+S�T�@5,�������}"���%<,c���&x�<M�����r�g�p1`I��&�)Ln��&Ҫ�Ԑ��۳F��o$K���&z2�}������f�
(%7�H��*���$���<_ʺTZ��Ǥ�k��`���E�~�?<e&7O,��)���ԍ�4h����z*���A���U