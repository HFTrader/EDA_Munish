XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5U2J(�|���.e��t����Tm�y�٤��3�'�ţ�N�h��N���IH�T�0��.m|	%�b�[�T��6<7�D���HT���$�ۑ&ܯ�c�H8A����|eb���/:<����\{��6�)�w��� ��pO�F9����ļ9m���^�����m�y�3:���&����1Pj
UUp��j]����0K;���M�t��ۯ���ǂ����|�������D�C�ǞnK���4"hfl�{J��g&��!\	Si�Ea��(��,�ߋ=!SA�ҫ�k��9�ey��<��;�8Ov��b�B���������ߐ���5�M�pj>�Q'T&�A]�C�}��٢�d֮}��y:��N��	�B0�4���(B��}�_t+%!��l��e�����+����*G�o�J��S��xz�) ��s�G���HDߐ�Y��إ���z+*�2q輄�( �d[���S���Ҽ�:����|��\���^�5��dV���~w��~���6 �x�@�NN�������k))���Ǌu�/��[rV).f*s#��S���߹6<u/gݦ�%8���٫�O-�w�\P���(����g�T�����=D�|��ͽس��}��*�u��l)��)Q�B��,E��r��9�"ɫg#P?�.��0y����:�{��M_i[4��o���Vut��H�G�y�{�}��E�R
ğ}|Nf|Y����g�6L#R.��Ϡ��u�i%J�py#�Q+XlxVHYEB    1427     840���� ��.5�4����>v���A�F ���9���ClS$h�(�%�Ke����s�^�8�V2
�a�sV��O;n(�N5c/�Ǹ�!���bg��I�o��#B~�#�?����/�s+)�tʀ�`���Nh���^�D�`P�
jH��O㷇Z����ٟ��`��1g�����>���^Hoӡ�EU �]��V�l��#;aO�6w�%��@��
��U��Xr�#�E	z��Q�o�#��p0��nՍ�Y�<[��~��󨫳�lIc�V>GB���2�D��鄎kĐ�&a0��qYK���.ʛ�#?Iq�Q0&s'X�8�Z�z�������7|���z?6X|���F��R����~�� Z)�#�>��"�H�J��	�~n�	{8�fǼ\s�x�vN��u�$E�pk�,�a�"��-�FX&bm������.�]�E�;�c����ډ���UG�1O�Aa�Jj81��u�^��� ����w�Zu
M&P���wC�{2+��.#����,+���;�^�v�8mg�8 �SS���������?a+����Q𩏻������J��ך����� ����`��Q��oV�ִ���i�T� �ַZ�����(ִP��wTkq �(8�j�ǥ����R#H�j��PI/P\�KVA?���y����;�d@�G�(�=��m$�H��2��f7=���s�����b5��P�f���C�����$��L������Lk{��#�M�cGDf�և���r�xG��_�2����`Px��ձ��9���̰ nI�Vˮ��'x����-�(#��ţ����<l����>�C�4���_��
�7=Rn�lc����`�]���ZP>�����a�w����;���]/� �4���1��
HZ��yݳ>����s�D *�U�#�n��^k0!H�43s�,��M�����a���H��
�fUC��󳨴* 9�@�6г��U�gF����&şV��9���4{/�bJ��d��3��7Ȩy�(��;CK�c)N�Ř��	7�{�ZJ�X���|z����3(�|G������y��vbP���AR�C�ܔJ+F� �B���a�,/����5~���[%�D2dK9�\$N ���{��ɴ���Q� �!H�oi'�6��BzS-�>�0���$���'�p�����sz��{����G�|�S���*��2�&��Ĥ3LzW{R���	��a���T�X��R�GI�)��ϊ�r��� ^o-Zu�Y٭�M�b�oblM��=�&dY~��h^�x�Ch?_{�,��*E7ht��ɒ�,���>(�������l�P��t��iK�����Gʧ>�]�yb Z��iYj�����ݴ�js�5�6�$m�*2�G���wt0�r�C���>**���}�9����k�*���
�r���s��* ~��;�-!3��JƢ���V�z-K�P��O�n� `����$吂�n5��c�|�>m7A���I�<�2/����kV��ʲE�;�&�ߣ��a��܉���0.kтqz���W����H��"I�!�~T!AGg��]�=����С��I�i�p���Hؤ$.�'J�}�i�	V���8�P�!W�=w���5k/�kļ;&x����6�9Κ:���g �@�Pt7>I���w��p�eu#���f��3Ca�Z�wi�1���)=�d�7�f���`!C�>�M�	k����2Z"q\$��U��� `����A*��F�`ۆ$Թ�G�Ä>�zb<y�Bb���v��(��>��X�]3k�1�7^wɠ/5ҩ��cQ���N�PiCN1�E��wV!�݀���N*�L��$��7��?�,�'C�Pp8���6��F�!D���6;�b��WF�.�t$�{��")�r�w���O_!�*�Kޒ���&
Й�;'֛��<� \V]�X}7s�8sch�/?�P���'Õs�%p�{w�-�ݯ	�>8'�yn!�<0��rZ�K�Oo�o�:<0	�LL~.��DI<�<4�d.��u ڟ L������8�����F��8�2�+�+�Bg�#�