XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���=r������ьs�QL9�9�z4�4��0��)0�%(���_�<�z��aļi�b�J%����;N:��m>FR�a�D��׬EWp[�_��}:��䍇 [K"۴M��r���v9�n�Wna4�p�����Ҳ��W�e�kˊNF<������e'#*��SVF����Yǒ�2�g��j��6RD?��rWNVm~��e����B��,xfE��AU��nx��������
�~��.}�7u���.����:��dE��8���Wa戅j��D�;]zr�}W�'U��/]�� P�%��3��ol,�7I�<�-�'�D*�{E�g�������:�9ŋ4t�$���/!),�� �C'����e�A	Z �t��Y��,8w�e,�m�1����♪��fm�UC 8��Og����}�^���b�[�+��$~&4zHꬎ��0æԘ�)����jDK�ѳ��>T�b��5l��a�\Р"3N���A�R|9�!q�A�}�W�� �N�o�Y� }�N9�=e��96��u0ն���0�b�aSF���^2zJg~'�@�/�~7���_}:V��lz�|����ټ����D���������3{���\^@FQ�0�l}#�:o!(�����s���Y͛#���>'�l��O���N�at�6��y�5��Y�	n��
��We�AF;��ԿȒ$<5��t.Ȏ�[,�yX #�>}<�Ex����>_:9)�#���-���״bk6� �XlxVHYEB    77d6    16f0l�?ʍ�L��I��;V$hE�8`ʜ.F.]^đjS��0W$�"+p�_2;��*N�v���n�rP$,z1�l��K.a���
��z<�G�2L��`=��A(�R�z;���%�g��b����Wȍ�xX�0U��q6�Q;B'���do�?�m-�"2�]c5oL�4�w0r�R@���y\$/�����/G�6^�/9�S~�Q�EzN�v UG�9�hfD��U���E��?��I��1H��F.�m�f�H�oհ�/j��7ݯ�I؃�E�t�+�l�s��g�fZe�X=Jc��N]w��C����P��HKjG��ݧ9�a���u/[;k�?��t�vE8�7/�	��6��e<�kq�T�}˒��� u�oe	s�6��|���ÊB�Y�[��9G�i܋B�b���B��i�Ȝ&���'9�8\�?��d�x�۔C��mz���TX{~p��ys�j(���`�UT3���Q�`�s�-A
�I��p��	��>�>�?; �^?g��i�uf���P��/M-.��4>h=RԔ�5�i�r�:0��X��G��54����-�d��ˀ%��Y]di��ӛ��� ���Vms�`������\v_H��Wn���K{�M4P�םH�Un�p�o}5�؝�`M��јd�E���	ҋ;/a�qm�R��g���UE<��e�/f�~o1_��Dŉd�h�~�~�}�6֎=
�Jk�'.��, J"��֯����w�t���62f3�x� �Ɇ�/�i��e��p� >r�r's�R�=��7�z2��F%ޙ��Uخ>*�3&�����,3~N$��8����Y&�t�WF ]Moґ�/�a��YV�ӕX�� �2����gׄ<b�}B%��s�F#�4p��=W����rQK�A��5]�����?�-��&�v�i�<eUP�C�1��ixZd�uΟ!M�4�4�a0� �ʑᑓ���=ȏ,̗'J�f�j2ܖ|c/T���p���y��rc~ ��'�������@�xg+ύR�x��|��S����c��ۢ���d����O����܋c�=��=�0�{KGa����"x�w�Y;�O�j$P�a�J��D;I�>M��6��>V�v^�s��!hYͶ�z0���t5�3Q٨��)�q����<QZw��@�K̳�F#g5A�*����y��奚�jS��O'���;�
��k!r�|�t����ɬ_�\�	��X0B��!vR�_�������r�?�#b�X��C�g~)���׸e�A����o���ә���3����l�H�q���<��`����A	��-H�<,<�Ӿ�ßUl�=��׆G�4>��!��� ��p+��:\*��ε�1NP�ֵ����@�+&f�/[g����e�A:��R3��621ik�7����U��*P߅����+i�&�@T�;�TK%,�pB�2O���.S��R} �NMnL�D�������X�&�Z0=%,�˖C�e�B�D3�ʡ�@��j�5(Ű7؟Y ����M�߂����<O�!/��Vϳ�#�'�$�!��5�nE#���~��a:�=�#������I)4�z��N�_�-�=c���!r���tnT'~)G�i��	q%~}�r��yl�h�l2�_t������^bť�i{��ئ�#x�cT�U�'� %e[���夃<H0=RVOp2T��^�F���O�w�km�)��y}��ԟ��󾌸���
���J����b6\1ܶ�<wbΧ������͖f: /Z��EѸ4	?9�R+8[h�|�5��{I��II}v�G�0�đh��~d�VJ�9�5��$Tr?�@��f�K×Dn�`�'=�.B�P܆r��'�W�,�����\���۲���ھRV
zbu�h9ڭY#a��KzF�#$n$Bq�|T���Z�e����O�J�[l��iCbߥ;� ��g�Ţ�{j;�`�:�JE������	g`� �[#��#`��R^&�c�T#ĉV�,}�cY�|�>�Z��)e��̣>d�E��0���^]W�/2��Ɛ�}�B��|&�h2�F�;/\%F�yl�Yǉ�yCʢ��z�Ҳ/5�v��X�����6�M����?E�~&J{|��dֱ9zPl6�8��H��5z�K)3j�YmZ���Y�i�f�]>?�x�-���HR&��є�x���#�S��^P�Z�ן!�;z���;�Lz��Ð������S��م� 7�����rq,�uB+Y˦�����F	"=����y%P(H^=�g�"�.�x�Br9;p������q�����`D]�%�[]�ֱx���qZ a��PČ�ƙ��^h��	B.a�)!����&������c.�Dl.,���ˡ+5٘��p49�w�t47}�[rҪ&F�vZb��	�2��E���4�g�}\v)_x�Ts��>�O<��2����!���+_o�P1z����[�߄�
��9��0y�v�DQ5:6�a?�=����W! �	�<q׋&sH��h��"}���6�פP�D)�^���� g"����ψclݪ�G���D��y� !��3#�Hć�C��*�_i��ᱫC�zG!�[L��F�uDF~�s����ֳ�˝�OY���i�2�m�����
��
w9b�:
���}g��������R�`����4N�ԇ�a�i��J��x�x;�<R�:�:	:�0�#�a�Bl��6
n���:5~�|*��d.��ܘ���.�KWΎH_:Ǚ��m�Q�7�V2Pճ�Xm?����3�����R@HӔ�h�:B��$mv1q�A}˻��aH�7h�)U(@iJO���e+�_�Sq��a�V�*!�"/� 
D�7�X�ǿ��8Z�u@0͇�*"���f ���9�-�@�
Q�_6��ul�����)REA�����Y n�R�w�;�+����Ew5a�8�Ҫ}��<*G	����!���[���(�G�u:�1���8�W���7�G�t�4�3e`c���@b!�>�X�͇A	�1b��~�:>s)9�����6�1'WɁ�( i�n�{�f}w���k+�=��:�2��1r�0ϓ�� ��-�4���[r�dn�@>��}A����-Ϣlv�|䔩��Y.sU�
���(�Fy3s��^X�n�v����^�f~��i�oǊ�tʃ��~�	fg��xϩ(��~d�hºِS0�O�<�#ܗ7�v�,��Dp@�s�Pom�n��gi��9��5&y�F���s��*Ulܞ�!�55_^A����Yp��@p��K��5&,�6�Z��NDҫ]�����ބ�1�?j�pf���{�0�]��e�L�B����}��֍c;tE)g�IR���t�F��O�J�c���﹓t��G��ɷ�YA�FO�lw����_{��Y��(�\��n��r��n~������:$���)�ڒ��[���i:�L^yiԀZf������W4傜��G�l�#�-�y������������rD�������84
ß�PC��>� ��z��l襘�@����ږ|F���f:���DOغ�b�&��Q�����s?�� ����%7$��o�)����I���&�P�S0,#^��"���:+pڮ 9�q-�LD"v;�"�:���-\�󔒅c�hL�yo>O��	�I��3�M:��X�nO6�{HZiC|�,LO�Ҹal�@�c=WƎyəo�[!uR@/G�`��rS��0���+���]M>�i(�cLc�J��_���)H5��[W�!ژ,�a�0A[�1���i���e��e�-o���[wP��/���B2���QǴ^��5N�"�Ӧr� \�u�0w$G'��"�|{�[�,f=����D3Û9�W��gZ˼z�螠�09Iߓb8�r��ln]pҽ+��-�b/
 ���9�^��������Ԓ.`·���\.��*QOq�5��?H������i�WǗ��_4m��^���z�N���D��R�x�q9H�����������{���-F�Լ\4R-8Z�j��-bo��H�1��"	�_W���.�����>�K9Z�(v� ��<��م$п���}Yy_v-k�5��!�H�0�P˶*��^�%n�8E��ڞ�G�.Z*$��g܌%9 ~��R�V�(��}�6$�
-[~B�T�F)��݄���S��Em����r.?�D�Y����9ΝΈ 	&ڦ�6c_��Wr������i_�~�y�&hG"���P�	ҽ�mq���r���Z|��/d�� ��3MA�_�Rh���}�p��gdZ�y���K@'c$gXp����A�Hѯ��(���ֺ�޸N�ӆؚO~�54R}�#D�4[���(p�uچ���������&�%���������B�f�>��t���.K=g]����ȋ�;�?Frt��8�
!
%�KrN\*~���Z
4����JɐU~�GŞ|k��$��+��N�G�9�'ݗ$P��V�������F�ei�;�?���`ox�l��X)fi���o��4A�5ҨW�5M���b!Ҧ����N��5?�͟B��$�N�#�f�h�G�,�o��n��zs"�$o���,�YP��.\G�b�R���S��F����s�c�-�@V��xh�r��)Q;P.u�b;�c�Kn�2�?�6,S��q���:���_�r�6�0�u3���5y�s���FIs�?��M�,�23We
x:��Dl��˘s
g�[^����/)��.#�|�;���,���_�AV�L'e����X��z��eKO���.-�]�,��q�0����ɳ>�ľj��C6LI�sgd�Q� �`ڙfo��+��O�ԛjav%���0�V25m��D���2��4�����w�%������+�����)�8��X���W����1�i���#ZMI�`7���E��ϙ2��V�q�����$�<��?,�����@ff	F-��[5�����?��s�D���eӻl��ު��� ����sգζQI����L"0䲸�N�X�����΍/z��-!t�z�,	��$'�q������(���:p���-��I��p��s��knsO棾㞼��p��>��&�h-��
>�٭���;�UP�	���x��1#�4�F� ���E�$-l����ih�q�'qi�w����9�^wx�'�K�h�Ub r�fߍ�B�
���@��r⒏G�}$�����s/#1{	��N���>��ȳ���$k5)`9ϨZ
�{����n�C�-Ueι��]y�@:�4��ÆjI�Ƒ��=���*�B�ߧ����DQ��k��@ks���f"���m=�@��y���������(���p�M�1Z���l{�4!��.[0��x
� Y�x�2bbbuc�+��mc[V=��e�
5�O�e�d
�k�7�yl����]8�C
�ǯ-/p�Y��y�WĽ�Ϯqn!�)ijs��S��efM�Y��j�qӶ�
��k�O���H��0j�I��+ɡD�u�|�͟�lχQ�&=�d�m��+K.{���hD \��~�f���I����׺�OX��xCID�o+�W����k�y�����mj�? 	��KiI�
����j�d�x�$7����P�m����w�KsB���]w��p;�)q���O�P�:>�jfT�%𥙙 wI�;��u��Sܭ�{~�7b�f[��I>4��P�i
��Km��tD�(�ŧ�^�1�E���rNzum�>y�