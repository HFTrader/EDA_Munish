XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ϯ"����պD�����5�k.�>�7�-Bj��y�5�OؑP���¶Y�����yܮvwu�k��tJ|�"�ߵ��1�� �>����Q���#D�k��X�\� 詉�f&$3�ѵf�� ��~Y�鏾�����K��Y���Ǧ.͒Z%�8��6���n��?�T�a�f���Tl�,��@@s�?�@�+tJ�Y(�m��RZ�v�����ˌ ݿ�S%gtT�*1&�0���c*
ʬ���D���ρ�-a<����R5�:Su�&ZQ�u4����1D`.�<�����b�4��V���
��5t0@@��JY�98n���8�V ��|Q�ǅ�%����l� �w��7.��%8���]m�$Z�Q��3��O�����R�,�[ЈLO-�ɯ���%�wQ��:@��"-�C����7��M�Q#�I1x0��:
��Кy\2�%0|²�WL���Rw��u5�Z4�+�SBI���;��,�ՠ��F%�s�eZA�kv��"�俞��SApz��4���H&�'��+h�pm*&���I��.�آc.iֵk����ò��5`�Y��y�N�hq��S���B=ktKXZ��"�E�����UWh�zE���Y����5'k׬�V~�����j
�{����=�-piu�tG�Ba
�<*�~���0b�}��� � �r��!ٳ�<��8��s�_�C�˹��DT	�α�xA�"E!n���W&�O3�_�i�n*�cM{n[_�-Nm\��{X�J��? �����XlxVHYEB    3d61     ed0QPaW��s��l����Wl����%D��s(u	k�sj�B��v�w��0��b6�ڻ!���%%�Xk<
���h��G_� ]����D')�o�oB �i�XYt��i���@����*n�yI�?���ob�@[&D��126�T*�-�� m�E>��T�������fF�-i�yx�g|�M�0�̂\��"��q�"[���#�3�JӲ���#��I�uh�:wBw��T�dH��1N^g͹�L;dA�l_����#vG��6�(��F�%�%��c��	�@�\��^m�X����%Xa�I�NI�+;ᄍ7i��N��K7�`���V?�����$ќu����l�%	�`O���50��`���m���QHF���b�������ǃ�be$?�h�p��~�k�̯��볏_L�\�B�/��QP��<�>��w�W�X��NN��+3�[^ ��Tɟ�ݩ��3Oy:�W��[Z9�3�t��1����0.�0��#������ML_�FDP���k��O��KQ'H]Gw�.@��,�~��� #%�V����1Pd��og5��ė�p����J��u��.&Yu�|�kD�5��o���Y�z�fpd���hO���j����>&o����8T����ƽ���	M-W��`���J���#�U:7����I���D)�y�
�e���!�Ǭ7ݻ�(�	��EݛgJ62v���]S�1�6Ѕ��1}����G�%q�Wa���LgF.#�dCdLwl#&)�J������cv[[�J_-Q����7�����F��|a�t������-g�Q ������7o���WhW��8At�?�����g���B����������G�j6&�����@ʈ�j���7ʞQ���m���B�yz�B��e�C��#S�N�]6nVߨ�Xv�*"jH��U����D-�7*�����eD N�Xg���� �����eg�C���4�u�we�8�3�ƚCቀ�3�;"�\^b0��^7��(��s\�(����%+�=d��s���T�P.�Y`�w��=*��+��F|�S�����{ͽ����3��ܤ�޴�[7�nÌ�G&��K�4e���A?+��h�|"�K۳�=90u�T��+AՁI��I�*�M�yL��
w����n��s�n������>��Y��k�9{*J�	�@ٝ�ߦ�泍�'@�D$"�oY^��߰�A?������	iw�����۾V��9uJ[�0�Z)� ��1�>��HjKX�X�q/�6~t�%}����-X5�Ƨ���@���h�$9b?�Zu":Y7�}j�uy:�w��l������+j����ޫ�&��0b�5ʹ�c<wa3�<�M�03�Ȼ�������T2\N�~L��7��I��U4n��e��`�7SB����w����9��E{`�- 	t���PD�� �z�Xe�Z���Y�~��3�r��_���z&�A|��

޵�0~{�}�d�jG�������Q�������	��i�s�L�֠S�h^^��M���:n���]'�fZ��2�G��$���O/w�q×<	7��j�oN`E\)�^ۘ$=z"����Ӕ`�i�z�@�]C=
�����Y1���W��a���c�pb6$9|��u�f���%w���?�o R�[T��n�'�>���4���������z��Q�,�G����D�����>Q<K�f ���&�D���0Q�S���83GMZ���A\���h������T�v#���m�=]-_P
��E���k�%��hm�F�߈N�?#�q2à�r���5�[��2/ơtD�~�*�5�($Gu�0�'�4�a�g/�>6���ǟ��;mfv{-�*�*�O�-�hPb�Ɋ��j����$c�k�W^��{�
;�������HcA�0
���_C�u6y�/}���	�{O�䁙t�{._~d۠��Ħ���t���y�i��na�ӻ���l��O40��s���*D��V��O���q�\[[���6Uy�sf0�6kTv�"����V�,Yd3ǒ�}��~2�q4Hͦ[I�g��2�1���?��N�U6ݖ,yO��KZ�'��h�Lj }٣�9M<]<�++��ʒ�5(t(�ȡٸ�#�����E"�T���2]k��fl�����4�Q]�j|�!��׎&b��8z�Y�ǆ���«�%9�m������,�oe� ���^���M�-t�4pF���ͷ�E���ۺW<6XRf�Ħ8^��4�Y���ѿoN��ᴤ+I!��I�<��)ʓUF_��:�GbE��+S �v�D�D˖O��-Ѷ���x)��v	I�W���͋}]y�gz\����"I���_T:�u)�o����9��.G��}��Ԫ���"6;t]����"�ͣY{'� CM �<ڤWGX�w,/+{��h�;XEB���R'zfk|I�6��B�J�9�j���M�����u��E��W7�����7�G���e]QֿCW�������4~� �'��E�[�m���w��I#;(8���v�0��M��ʟ^=�'�DQ1UC]��v�9�ա:� B��.��� �xU&�HR�r,5h�֡6)lu+��e�k�<к�p�zH�.��~����>Ȣ�a�=y�ca�7O�P������8��-��(�6L�{M�#!��:����t�I5҃���Ǐz;ϫBE��d����N�H�hRҚ�2���ʵ;� ��:6ܠ@^6�B>��)z����Z��p!����S��*n�����L(Y?5�r�S�EPsO4�����4��&e��d�J�47|�!N9:O� �f��q���U������sDs���g=��C�-M'c�j^��1D�$�i��)�C+늎�b�w�Rn���H����R�4�.��g���,�΃@ -��Uޡ�`>�xAJ����Y�mn����A��mω[�eѠh�D�Ԟ�y�7�F<DYx�t����yQ9�� �H 	G۪���x;�P4|�a��iE�S����@"�W�G�#��C�~��m"ݓc�>*��嶹����E�ǝ���ؤ�Cu�N1�`�B�����:�9����G���e2�LZ�b�chH�ht��u��S��1�*4[)�_�[w���:�7E�@8����k����@q��KX9R_so4���:fjFlij)ڜ����4J=[&}}��.��d�1lNk�|��Sǩc�^����@U5��1�a� �=�:]N��,Z{ө �̦*j��jjfJi% �҉{�y�"�g9y��c%N�q�"��{��6Qr`���(��U��TC�=.^�~?tsB?�x�;և�uM`��;���"UT��y������{��)�\���8!:e��ND��٦�������wjӞ� ��@
G��c�g�5���(Ͻ���&�P9��{�L��SĦ�e�Y� muT�Ũ7��QX�K���/ ��ϫX!rl�u�ȊU�/�x�BR�0�w�iA۳��N'�0�#q/7�̘e<&qIWX����[��"� ��2�aAr�ECǾ�%���?�vP���)x/4q��æ����r�V�����k=L��[�G���3}J!��ᜲ��w�۞;��e58x��_R�ҭbGm�DZP�{ub��������O�����s\d�?�O՟׸