XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��xE�j�)�\��z�:
XB@9L�2#��C����j\��S�x���fs#�?�7�1{��7Ff7�����t4�wTY×M����ү����ISa�9�>�8MOȤgzت&��q�V����f��b�F�/����eΊ�2����-z5P�]U��Wm
�� �%�w�s9`O�����D�I����A��8�['iAe���̖G��I=޷k��(n�=����>���p�t����.c��&���Xi����zN�2�Z�F�<��+x]��|����U�B*2�զ�a�)���O0���U��cW�U�0L�.�)���А��Q*�^ֺ&6;��@4�U� �3u�l3VD� ��t�� h��laI��� ���v�ځ�E�7�t[ґ�Xk�&�
��Kx5�X�LP�Y#F����/�����R*}
��k�5��b-̵���㮌�5s:Ä���j�siY�� ���>΁�Ì���a�K{�Ӎ��'/��0�?�3f�s�-o��⸌��b�@	g�;�D�-d@�?SN���7�J�	p<�Ǧ�[�?KVЂ�Ь'�dNq��;]��sxע�6��/��ٕ�%���?����3�	3��Gf�ΑQ\Ǩ�=�-+��\>�A�J��O��z�^�LV�5�8�ݍ������S�TD	�RB"�럅���:$p�+���z.o����%�ty�E�$�͟�P�EەEx6 pM�"��T�B�{P��GJ�&���~
�tg��{�"��Y�fŮ��	;�XlxVHYEB    c3e8    1d20h[0��	X[��;3��aXaK�C̡_?�fݱ��-`M;���L%ʘ�~�15������Π�ů�"d��Fի:��D.��<ƿ�[ڏC� �>�~:�[��u5C�3��'�ż�kP�\��Y4����j��z��:��KH�o�8�2�������{��%M���[���G�VI��x��#Tbe9sb�J�i��iBo�yzt>n����N��?f�������}m[\x��h�h�!)0������$q�-� ��IK��)f-����V��L׮e����d�a2o`A�QBU��R7`��x������E��� �P���s���`��dЉ�SDZn��l�ע�ޥq��p| �<��폯��D0�ʗ�[hő`��j�L�Ҋ�ga���A{M�b����fi���+�z�҅���Yn]�bh$g5�Vo����Pzܓ�͋�ÁG��w�����$]��\��]������l8p�7�O[ɨV��
6���jC���_�^��{����]��˗�V <z*�	�:�zk��T�����%��c�U,XC)��n�C�ג�z�	��QQ���;�RIAf��� ��Us�+�oES������(n�߲���P�~�=������>9UЋn�����7��^��cV���M��e?�%&G_j5{�|�w Yd�ޞ�3&�'��I$pc4r�ph5�FGF�/�>��{�5AƔ��@ ��!���4S����*�;Qho-J�4���ԇ�����4�5�++[�1�$t�+DAy*}�8�m�M��2�êV	~U����7q4���M�X���כ[m�0�ӇP3��a}L)~�ó堙QeLą��B�%��T��O�LJb�ZI)��پ��Y�[���Y�ʒf�	�Si���A��Ĕ��V��% �*Z! ��w�k�)(�#�8�+@�I꟧�cr�>�������ڿ���gԜQjP�gP��o��=s�&�E�44+�M�<���~��wT�ꗁנ)������RЏ�x�� >����F�Ayj��yռ�V!�W<	W��8(z�m�s{���V7b6ā�	E"A�����l ��>��@,�K�ۂJ(i��%I��9jiG߳����,�X���Y�zcp.U;Ǟ��N��LN�5vڣ��s݇4�����9'd�,�S酪���RKI��u�P� �A��s7`k�iB�hsH8���h�R�S���ՍyP�[~�<�4���?��q�.�M�8�\�xhS�?��YV�Qcu�1^	{�;3TnAI	D�"m��E�ȝ�by�����m|��S�r4$�r�Ζ��z���`h��_bmH֋�{u�R��T2��
����+e��m9R�~5�Vݢл(�hr���j�&U�Я)��q9hd��;E�ט������t0Pt�e^<a������=��k�.x��qǃB.�E÷�΀m�  r�`G
�(Q�_*���)��a�[�Ǝ><�婖�\[�<�LazC�> �� 6c"�R;
����t#�N�����mj�{�:SN���I$c*Y���JV�/+2���)V�ab�C�k�=��4x�λ�e�C�F�<�B�Ψ2�G�08/u� �����K�ܮ��F~�E�Z��˝1�!#�!�=�w�U���n�ڼ���)2n�貊����d�e[��4m�Z�yi�/�7�	��T#>A�jǊ�l��AO��0�_�/�wc��MNWO��ӯ�[x�2�4�p��uK�H��|m�r�M	�,��f�����u�4�I�y���T��_9�eKF��qM�{z��Zl�ݏư�П��`��Y:3�f�q��sf���G��D�"�n����q�|��U�ɒ��0�o�{�49=�C�{W�D9̍/]r��	�Ȃ��q}X���`�x�����-�q�����?z]#	X� ��q����~P'�cIUn5� ���[��0hw8l� �Ȝ��阿��O_7w�}}P1�Z��;�_�/%X�3#E�A{>�cH,���e�׿QP�Q��kmV�g4���d�5���!�����h�B���SiƊOn�ц�`��u%b?J/Uڤ0�P�܌ V	(�F/;�^�<���y-M�)��Z�#��8����Y"�$�j��w~�}x�L8�\��t)%6�(�����/�q�o|��C6*�~*.7�;����RK�f�x�/�/�[@��P���P������7�\�`�[`��"��A�εd��~߿��̞�m�"�[
�S*�<��`F���f�k�꤆�^��A����rg?�+B҇�'�N���WC3��xC���I�w�sD�s0����!(=����{Ĺ�%a�Pfi���.g0P9��F��)%�2v�;M�^����+�6�6��/�B�cr��=�$u]��N!�d$�Ix�2	0~�6	�?��,���G�G�r}�b�aPwaN��=O:N�D�%^69��T���G6���Ft&�I��,����	67V�;?����#�[���~~�n������Y5���y��v�|v��^G�����cRT7�#�f�BH7��U��-6���wF<gJ!-�$���l0m߂����Sk7}=��l;�}X���=�d=��y��*	���r�vV\���L���;���/zr���ö'����Ɉ�Ŀ��}y(W[�a��?Kp�8U[7�5�۟��$vԝ\�4��7sT��ƲD�$[�k�^���>�_"&�fo��I�t���m@3��5��n��`b�/�q��gD&�P.u�0�0.�JQӫ����>:E{��,���� Ų����ȕK�����Łk�<�|�x��	v"ґ�|�z��&z(�j�����h�k��j�C,H�c�PR7���A|��t�N�j��R�C�@�0յW���N�~,g q�V�(�!7��_7B�ѥt�����+1���W�������\�^^�
U��,l屶Y6���(Ӊ� Hl�(�>�-��CC������M
C*$��v�\�I0�t�eخ8��|�����~�����9�V�w�A�s�X��~�X{D�@)�q��\�^,�>�0�`hj)�&�Ј��K�Xy�K�+]a��2_��2;���'k�z $g��R<���b��I|#G�����VU��H�v�k��\����(b̚z�"�p%!y�<\I��j陶�l��H2��[���u.�=�Ě����POh�D�Ƚӕ(�HIM��C���=ܫ��b�I�s��Y�狒�)�=,�{@zoj�4�ԩ�����T��_.��ɜ�/��?i���KӢ���o��xLޡĖ�LF�YY% 4�N��D?���y��d`�^�X
UUّ��ɢ��gN�b1᮷B�1�<���u�����t���HyQ��V!S���<��V6����?G�
�n�|_)���� y�4t�l3E;vD5�?_���V����Ҭ
�W�j�j�i�Yߝ�~b�%m����%.�b���%�����|��;-I�˼�����H	���t�>�Bh{6W�%�w�����\�'$������Q��>���P ����)�jw��PM&��ɡ�q��lDE�s^��3RMe��\Ӿ�?2x� w���AN�0�l=ԴR:��á�FU�'�u�. �N���<�	P\�ڔڡdD���8��׳�V�{�٥Q1*�)�o���7��K��X��a������Q�"Ǫh��Xf�S/��\��������X����&~�Ԡ�(�x 2���H������S�3]Ŝ�������͋<@�ѓ��ޤ\��c�j�Y��੷���Z� /��!h��������Gt�b'ik�㍅��-��^G9Ѹ΃�haS����Ze�`������=r��������9,b{�[U�h+�˞"�"�f��z�@չ�,%Et�a�l+�ؔP�{_�nO=�v���3`s�ى�,�������{�HfE7�U��gL�����:�D�>���:R����k���B�`I�����)ӹ�P�_t�Ą�`T��76���rYG�C�U�4xW=2>���hܸ9�t�0B#5�ӫ�V�p�zJ��z�s�' �Aܧ$��&�C������=譽v��zͭb��$*��Wܽ(��ѦB��n�e)
�mU�ڟ��iI,��^q�6��c�lΟ	��*~,���k�1�d&����{�?pG0�x�[�i�pq��Я2%ͬQ�a�K$��O��kש
�,Q|h�u�}Mb���WkY�f��aa�!�(�����ϊ�U`��	��J��Э�*����xDGC����(���!J�s�^xbW�L�׳e$�0�whF5|���;CD�����_9��m���{3�*��4KJ�sQG�r���z��B۲5��KPO�^.��Y�Y1��w~����9,�N=N@#�y��1�R�7���䗯��.MF^�,��aiR0�"R�n|�/k�� �Y������uÔ�[/#�ɻ�MQ,E6����$�Js�̛���^��3v�u{�m�©�t��Q�pE��k �������i2�'����F{�� ��}�&Z��|��@w��ؔi�η�~�0p'P��aH�]1���;8�=����U���� �#�R<
c�]��e�o6Q��O��9\M�$�7��TߞM�,�ngm�`�U3���(���FL�jI�~9���y��.f�|�(9$���wE�j�x��fCD�l�4C	��2�2�ي�fVĽ��.>�o��9¡�K���i��9EE.WD
<hhZ��$]=�D����1'�e��,>ണ���MO�5,�~D-��ﬖ�D���go� �\W#�T4��\c8��eA$��N$r�C1e�k�d� �T�є�D�{ph+У��iA�ֻ�6�X5\��8;%����Pd����{�����!n?��Q���������@�H���i�:G�V�[��^g:���`���ݵ��b�TC�4�]C�����\B�޹��������Ȕ�+�-��&v%�e��yN��_����W?)�.A�=�3�+�Oo��];7)�w?3��@��R���<^�^�t�AK�ߚEjEO��tؠd���(u�?=���������@��ۮ��aCrd�&b= �#��Gǘ��I�s~���}��<��q��*yD����C�������M�sh��y��c�G�?ΡӡC�������J�S��$˹�jU��m����y��%'��-(�_��RC���n�̏-`Pf�(c�Ds�g3�|�A���grx���3��� r��6Ӑ���x�ɼra%�<���yk�O�����)��cR�A{��6K�.p������
�x��I�#IOQ�*ֺJ��m�I[��U25y�����*Q�q�J����� �������f/��g��LF�W�CB����Ǒ�f���?�q
�����Ё��M������p�0�By�����1Y{�B9«4q���i��A=U����;� h-A<����v�5~&VV�B���Vi/tWb]p]Q�v8�ca�sdOk���P�a\ r�������gԄ�e��.�g�����.�c|��KC0
5�}�)
�ifS1ݩx��R~6���!;�$K'.�y棸8���T��c!6o�u�%4���Yv�ߢ�J�p��.��W�Ό�y�5pD8�Ք�q<'�sQ˘{&Za�{�����7��L3�pO���G����rUj��|ĝ���M�O/���n�+�D�솓�iwn�z�И�ԬkG���L��I�r����)q�J^l�!:4����p��~e�Y!U��TS
��_��#oΐh#�A��䆠�D����G����Q��z�l��8�ZoLP¸�x�N��e�ZO���"g��7�1t�8u�� �^:R/ri3C"��b��T|1��k/��'��k���>}�>o@�8k	��n�HR	��^ l]�+,�D�G��.�0M��� #���Y@��7ث�M�kޅ��;k~:��W�Բ|`d�� ׋�0�X1�����6����8�1���BM�;/XB��&�`nE+���a6��y��QͿߥ�Ug��[y� �cH�)_.h _�)3t$q����������n3��=��!���
HU���X��i�AvBc�_�҉�w�%	+u�w>��e���M�-j��%>��d_N0��������S���xP��ӌ�2���4tl�%�����{����P-R������6�.h�o۾��������4J��M�e�/���r�9�'���LLV��ݓ����F2��y����$}����F�|���!�/;�������z6W�H�H8���~��)zօf�1� ��3_���l�՘0���ɖ!��cl ֶJO���"��7|���ԣ��4�^v�2%�TUX�ȕ��:B�S��wQ��`�
�0��;& I׳�	]��?S6G�F,0���딋�$��]R��^ziQ��H)�T����'�����0��U�To"GFF}ڧ������q@sL�E�U�F�*���B3@�o��	A*S�{p,`xyN8f燕�BB����d@~�7�C�U3�������0��vWp|E���̹�94-
��x���x5�w��k{ǹ
2&���-�L�?o����f���i���t%�}���|_��s����Eͥ�!V����
�v��%�,9�e�.�	^�����P�&�fX�I��b�kmɰ�f�rR�R>P��U�e��6u,e���Vr�}�]m9��3��IA|	�'p������n� ���(����g�!͂vu��25W�ɫ�O�Wo]^P���d���HJ�����W���n
 R�-&���:|��v+����ym�G�0T���w�߾iѾ��<��[#J�0��Ç�P�<�0��	ԏV������i��M�E��BI}߻:��]aZ�a��K巕�\*�7�kGU.�}\H���4ɘ�A���aX�����T}�>ۉ��2'�Lj�w�e�9��1>dF��دj�_�ڎYNGr����=U���*!2X�-�eBU_U��[�#u�?����8C�Ϯ��v�����`�ǧ�H�F����Ħ��&j���0�r�t�^�lE��˗vNJن{����V+�߯˲PZ�hÎz�#�>��(�E�N&�,b���*�
ڥ�z����P�}���|%� %o�R�L���#��;�.ǧ��U��'-e�\P�Ѻ����u�5ᴲa0��;ty��~R���C�d�J�