XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���U�82�ԕZ"��s��Vu�'��*�O$�Z�HQ��>lQ]h��.t�^������ʑ�o�2�/��o^u\pp��=mb3��7��03�aA��D�o�	Z[kNEQ�����8vj�i9Dq[�:)O�rH��@4�#�z�qC�G���Q7����yJ����a&�`m�!�=�J{l�M�(�P�l�L��7=	{CL�Y����/@�Vϝ�Rf*������V�GU��/�Þ5��!�-���s�^��`h_x��2F4r��G]��:��:��DWTf���Vwp�^kx�%%f�]M�r=��ݬ4��;:D=����F����z4��T�+��cH.�d&�&+��F�f�h<���V]}�{a*���S�Yal=N�_�r=M@
�JÀ"{Y�U�۠��(e���EZ����L�~fAB���J�lo3I<�m�$RÊֿ6e�y���9/��`݌}iXX(�M�]��17b��Pb5iw5:�4{=��Tھ4��488� _'@���L�X�J�ְ�c�J�Aӟ'F+e�em��*f��7��wn56>@�;+�3�����zia��ܒ�v	�ST���~��<��u��	��l��)?�fe+�R�|�c�^-��פHN �v�:	�B����Lj'��p:{U�]r���N0�b'�~�lğ��3Z�hG���N���ĕ
�;��|�������_�4V��Ͻ.&K1�}����C��L�m J�wF��m�W+��Js7�◺�T+�̸��2M�XlxVHYEB    fa00    2240[�>���2A�2��ɑ'=���~�픣H��f�2�Rو�~��zB�������c�)̝�K��k
P��{	���z���(�>9���"��\�Rl����#��&�<`۟�T�Jqn�p!�=���FK�k�~�
8Nu��E���_�~�A�b��mJK-#��
�I�f7�C��k�8�!�jPs�5֣s�m59�j3�qoȩ�v(uU������i�����ි1��|>��h2�"��U2�* ��F�fh�%�BR�%�2P9�����G��aV�T�����ҹ��jF�#����6�.}yq��aV:_�:�y��H��Uy�K{�W5븬9���L�u/��Q��ݘ}�I�	��&��#$�щ��_�l�[�K,����W�4_�����G����ۆTϬ�Ύ{�g��G�P��m��`J�����.gFNUڅ�q��
�R���e�ǋҏƷ΅�տ$4	}�O�Q{)S��M:T���~�iO^,�~��<;2�n5�KD�F���Ұ=ژ!Z
�`�5��x�پ��L3i�U+k3���R;B1;#����O��ȫ%o]���O��`#3/m.�Q/ć�%OQ���xxذk-�Av�֛�5C2Ex�������-�6��<��sʸ�������5B�	�A����Sͅ]X�^�Ѭ�<�ںs0LR�N�C�=*nz ^�;IEBX���%���V�1cuW�w�:��1^i�"ۑj����J�
�Q��E�k�~�-+�ZKc���Ѐ�5��9y��BӀt��`F�x�r�hU�w1#G��(��P�O$�ab0Is����Q���x��&��`~ Y��9"�=Vu�גh!�F4N8~Б=I���V>m�m��|�x
�YZ��]G�#w?�_Z�T�0�rw���]�Bb�R�R[�vV
���V��v�w�����9�XS�(�*����Sĸ�h���?$o� �޴}K�~I��*��1̞%y�*A@l�����T�V�.猇~��!�����F:�A
�D g�1�2l7u�2��J�Q��<0Y�2�?��Td�n��Ǳ6�Ӧ����3Z�b��/��mt4P���.%@r�,s3'���غ1��?aRat�p�3��8%4#42�5����{��	�탊��c H�B��kzT5/knf�F��N�""�NC�y|�R���>X#�Y�p������7��@R"�����������bX��6\��ܽI�>#5�oК����f�q<Nu�)E8#��`&_����2�D-Q�t{�D>�����Qf�� ��3�p���aWSn�w'�v&��pE�)����(nnK�"(t��a�H9_�y��*�pu|JZ���7�7�ZI���~^!��7<%�Zfe&��l>��?�1�M0h�w���Ϛ։ ����kl3R�������G�.Q$3���Y��e�|o��w����B|�1�w�׽�O4�c/eS��ZvI��4��,��b�$�)E)��e�������"��΀��.QKڰ�m����㉢R��!�)le��⍴r|$��oUwD�	���8��0v�u��j�4���o�w��;rıI吱: ��	K�eR�KB5��I��~����ܵ���U����<�N��R����*i��Oc+N���`v�nC���|��=b���
'1��M�����Z��{$�!���_>_���p�3G���G`kn�B]��7�c�"�n=1���wxr�����ԇ4R��r s'9�q���_����W�FG!���=�������4Fl�R�M�Y�jaߛ:b���MdLvk��}j��kGW�ݍL%�q_����2ƈEs�G�~���V W�p;z��د��bR�eҦ�D�3`��!%�T4�(!�q[�v��>��t�*)9�Sµ���'�5�x2Hx]A�v�-G((VR�4I�d�ՕX��s��&��;L�m�E�@�C����I΂�pڮF�&��߈En�0�ʞ�����e�}�Xdi��0{��Z[g�K%���S����o�F8b]U�Z��Y*�Q20�2����*�b`�(	>ّ�՞a�Eѫ��J�� r�߲$S�\f=���r��|]�^..�@��
��=���]��O*Q���Y�s+�;������|����F�PNYVl
1 ��N�kRy�j��Yr��pv��a�}0U���*��n���L@��`tY�~��a��~%�{�~!���݌�c��t�>��Q���" ��ۂ��
j�)3���Գ�,|3�c0��Rr��1��k����mDq��y��`�GT�t7�hܛ\y�(Y�Ӯ�/��9`��H�]o0,�DP7�����yV58C4��݌��j�|���E[���W��v����$!�����7�C� x�����]���)�* ��<=�+����P�$O���">
@��m!8�<,t�	�e�ѐ�HC��c+-yh�����h�n���m���~�}������R���n��#����rgg���(�_��Qw��{ȈOo�	|\K��Iok�e�<Bt�1��<�7� U�=�M�����t�X�Pu�Iu��>%�Aw}��[]��MFS��Ɩ���X��д�d���- 
�fѝ��tiL��D{���\s�$r4u;�q��(V+���';���z�ǃ��^)�⽹�6�,�*k��fŻ�:W���^�ڟ_�L��t�3�Y�j�[Z�P�>v�Ͳ5�#���b��MC8/lԨ8����#�y~��
�[���>Î��(��99^@!׻c8{b
��j��<�9�b��҄�K�L�6���#�-Q��E����U(i�]-���4L�%F	�<���T��[dg%C����
�D)���{�Ɠ!�3�7%��^�M�����تƸ�(�J��Ճ�[��kԜ��l���9��`>�����ޤ1�~��$5O�v�y
qk�e���X�<��\ b�3|��Q��ݜ!��hYJ�3�8<�� ll�p��l!#��˻b����0����Q���wV�2�XS5��CE��P��\���:@�ǽ��%%��u2�L:*�^���^�-��E|��Vt���� �zm�4�h��Y�I@^�gIP��w�T�(x ^5��a��ĝ
�A��HE,r���[�A����N)�B����"ʳB;1y�0lk]�f�4 ����u�9� 3�G���1$1�֑���ٵej +��>)�Q�]��YփiZUR���w$�Q��Ÿ)<��g��{.��)WBh�S�$�C#"jj¹U'{Oʅ20z����K�^P��1��lԡ�xY�܉���յ��A��{�Oo񀠍Rr�7�ZY.f�l罵1Ҷ�k�BW0I�T��l�!Tۥ'F9�K|���Af��P;H�tu��n�:e#eI�}H%��]9c�!���+n���'��|�(���’�%��Xf!�l�+p񻻻�.2}p��������
�Ԯ�&A�>� �O�~�)z�;'�8�Ox'8XXZ�+�������^�.9o�����X��:�u�k��}ּ�VG�V��N�Q&z����JR]1�agey�����L�] ����|(�_޸J'�Z:D���"Cl}jo���KF@��� 4u��n�����\�e\�i�ۑާN�0�����X�RJ¨0�[����B4GEj�v)��D'�Q�T�$�8����czv��Y��֣�_���!8����-R.��u�B{�4�E�CxIAݱ:1��x7���]��0ho�)��쉬��Oݶ<����ɍ��1��n������9��og��p+j#��t8enҊ2đ��z/d$��d6ʸP�%s߇��(�"GzHcz��3: �_V��v�ܔ[�c]��>|5B�lo�&xm��O��ڞL��4�����G�{�Џ�V�18��{j��0�:��U����4(�M�~�/18g��I�&��鰼��<mn}>0�]Ys���}�)^I8�XaW�� ¦��a"�6��=��B��F�dS�n(�2�$�����9
O�O�����闈dĎ�͸9����%��I+�^(=���cQ�Ӡv�|�
h>>ñ���@�W��	��w����1H��k����~W�t�fb�B��ܹ��2���4�Ci�<
"��MsO��熟�2�9\�bn���j�JR�+8ʌ݆KM��%WmF�J�\aCb(��&!6�+�\�YW𭋼��ƒ�	�[YJ�VIKF����;��HtV�q2�9=�6�Z�co�sJ����X#D�Yzk�
^������h|�����0*VH���ެ��}��c�+Ndq9p��Gg�TP���r�2~D��)���y��H�<Ct�p�F
U�֗M�T��x���6��IZ1��Ӯq�U��H��'�W�W��ڮF��!ٺo����ku?���[+��l�{{�5n��~�����[�a"O|���b�Qv�2b,D�O�ٿ3c��
�1O"[-U�̫�!��.��g]��v�?-�J>�K:�3ͼ.	�{c�Z¡��8��x���{�l'���K씬#�ș�-��f��)��`*��1���1
B�V����E����4�x���.���R�ğec'^���?�
;V}7��0�uZ��!V�׏��I-v	R��3b6l��@O��	sZ{nKDȪu�Z�/K���>Wu1�Ȭ�D$�����q���K`Z4�'��Ͱ�vc�l�L0�)��|��Zť?j"+8���w�m�L�s�K���vEH�13LG�tG��meպ�oJ`���O���<6�e᬴�q��%����4�Z
X�|�o �e3����qrƩ/_b���s���ɞWVC�I�#0Z��yZ��p�ݟްt�In�{���D��C���n���E� ���BQ
���`R�M�.pޱ�Y��s��Ǎ�;ݦ�[x�0��{���"Ң�:U��ǥHݴ���z&k����H���pT��@{ b�n����.ߺ}���r���\��x���,�a��j�G� ��)�J�*l-��~R����?n��ͧ�j���^/�!j�{4�v\%�m��?'�UgR*"7����P�q�� ����L|ʎ0-D��ֵ�ڌ��X�dX����u�#ue�c��$��v�.�R�t �2��b;�34XR��c��?���&f��5�H��P�����)'d@B<���^m�����¸�Ç��vQG��K�ʷdR{C��槸��c�jj���-eF�b���!�t�],���I��v1k��>ɫ<���N���'�!J��^�!��|��1�l8J�.��\��J�b��]�_�-��6ؒ:~� /V���/�c�⩐?��!���'�� �P�cg�Hsj =Rϒ:*�mA̼dCqh�ܰ��:B7����&��0��gy�3�ؑ���#߃��e/�����Cۊ�H8#*�=�OS�Y��]���^��iάzK�^�B�.� �@��`�I�j�V��dU�G�%��p��/+�B?#H��BUHݻy5�>gB��*3@�߻�眰��^��Ch��]��cx)qC�;p�T%�m�L�tޛĹm�7��U�sS��wfH$���U!�]k �P��P6[�۸�kj����:/�6�����p	��o�HH��s����t�qd�Q�6��A+~��8N)�@��W ���h4r�����i�~���5�|��Ʋ����jb���p�D
�1�.����"蕍���Ӫl���o�V�k+86��&j� �i����ud������&6ZX�JVT����=�N�����)���~g���B��e��F���t'&[~��J��Ўc�־��tq�g����̼���wѵI\'V��t�Sa��uAvnE��MuK���D�>Q���C��'ۻJ6��z�.��
ؽ�&0|�Rϕ�8��Am3s'KM�A֟�B:��9F�K�� X_��p����F��f*f>h+Hd�҇� ��Y^��p�!���e,�[&� H�̸멞A`��X
N�j����"��d6�o��b?�t����cC<�{�h{� usa���'���Õ�!Ri�ĪuX{-��|��#^d=�דxv
��>�;"S��梞hP�l{��U�U���U%�).Q�u_�c�y�H���;B\��>#jJ����@�e��RQP:sK�tc��.QD_�t=Y�!�;rs��a�͝��޽�����XKg������柵��K@�! �A�q����2�#N,������"�Qך�W��\k�xP�q�Gj�WAM	/ᘍZ����RKz�yƟH􋓣��|]��<+�O����vw�?���H�R���&�{�o?�۹G�}��Ļ$�"3[M��V�C�)�Qоzk�՚?C4\�����#��y�����w2>[�lwq�Lh1���Tھ�C�:�yB�_5,=���";��3xQ�r���DvR-���A����H�9���3�f�W�����8_dd�[�?�;+6���D���2�x��H����lY�G�W2���w��缷�E��!KM�pm?���{[y�G��w���;�����|����G�ؐo�G[�L�i���-����ޑ0kC��yT0�n��#�C~��F�4�J	+t4H� �� �g�l=��� ������ ƥyN��S��*
a�I��H2�����MBFQ�a	��dT�$�*�������T����c�G�)W͸�|�V�^�ŧ��or?�DZ2i2����Di��\r앦>��O;�A05�m.�����<aK#N�B�.��20D�j����!��0h�+����;�|�|���\��v���Ui���y|��ٴ��h�7���wm"~1$%��^%�7X�r�̚F�{�P%'T/���}�5Z�Z����|^��"}��v�.���_K)4s�[�k >��T����}bʯ�P.�/��/.���Ǫ�*v64��P��.$��X���j3χ
f^�e5�_fƖ�D����C%v�����h�>)�����S�>���s�+�'ҚHbŃ�uG��:���2��(�&�s�	�%$G���el��ˌT�����U���m�Ѳ������{i��`I��!Ϻ+�x�3�����q)&@�D���@��ͭ�s�z'�e�Y�F��Q�Б8��������+��?'��ִ�o��킩�K[��<�䀰�UVU���r��5/ٌ$j�~�h��X�M7<��21����~.�fzf%��Sr�O���d3�a�.ͅ��*P�:VHz\%U�1���Rr��uE�\͂�͛������At�ܣ�2�"&��wf&Z~L�-w�{J҆�[��r�A�NS����9��5�M�B��/Tw]ώ�p���`K���8
��vBÛzd`yN�Q�.o�٪]��	�ִ�Ұ�ఌv	ZT'0�dHY� ?D2Q��z7�
��X����W�7,����b�`�Y��m��{l�Ԭ3�����^�q%�O~_A����C��|�#�C>��Sfb�˵���5��'U�����޶ ��f٬an������
$"7Q�<�,�p�,r���檥�-��h�w}���U���<���Et�Kd�/���,�I�/�r@�॓c>����C��Ƿ��2����^�
�|`L»N��6���_�Ya�ꡞm�,$3�M���v��<˥��&t������O~p����j�f!j3�ox�z��e�����!FY�"�#H�'Ka�eO9R�ܛw]3do��s�l�\`f)�I��m�����Y��͡�ϧR����#�q�|� ���U��A�;8S����}g����^_U�u,�sՈs��� *XB.t�/�c�P�FF�X'P�X���M�w��[8ڮ&�I���צ���E
��!�äf(�[s�$�
+lX6�V�� '��E~�zm��9��|�pl�64�U����u�Pe���5[-���)�t_�X�ƚ0�yC�+�;,��R�bazzD=f@�E b������벗�7��cPb�/�3|E~�#�q��ٸ��S���N4�|����lї����μp�r�@���͂ٵ5os��V;_�痲����+�'��0��f�O��u�(�Ս�ji]Z([����)�7�0Z%�%\�Q�8޾N���ٷ�qR��������=K����<c��U!!X����wf�4߿|����e�K��b�M�[�Ka:�:F�1�Dm���sz����˨�$4�����%��i�������!���-�����J+��px0V}��&�0��e����I8�/�����蜕�)����)@`�
+��l�I�/Ͷ�)Zfy�gO�m �Onu9�]�&ruDT� d4߽\��; �M]�hr�~��+���~f�E��v^u�x��
|ZǾ�ኼO@̉�/qƵd��izx|���� ���b�3��/	�ձ��(A��P����%�(-"�i�/�/� 2):	T|P�a�⼙|���ۈ]ў��be��%�7��MM^��J,�&�b4��Ae�-b�9N����ZXlxVHYEB    6682     5d0�
l'OY)1��詀n&�$���&�	/�C���A��E��O��l�_֯�	K؂41�&���|�������y�F�Rtm���i�|'�����%ݫŸ�x�=��,�^9(�q2E�/��=��ώ��[*���~�։���}���rV%�X��#	�=-˗j[.�P�P3�_�3�����D���+��F�-I	�1^���E���\����	���o)?��u¥d2B��.��VI���dǰ}6hX�F)x+`��9��~n%�zP牡�H계���('�e���34����8��Ts�!<vs��/D6�\�����,_�Aǵ7J3���^��1������Ƨ:XD�����V@�n'6N��Yw	hI�]k%����)�	�Vֿ�&٦�o��5w���V�6�I�¿@�%�wP����'�"{��	�@���I�Z#�?X%�װ������rʖ\kM�0�����e����@� �Y�
���.z���
;A��$��^�5�/~}_\38t|��*�Y�cRV�&o]�e߹b�%Ӽ�����.�C��L��s���Lq� 0r�=1��a���Z��]oT���+�SAU_��$�$��\�C�lh_yD��9�l�WKw��˶vݿA�P�҅aI�N�^7c^;S�X���|e��o*�|�O�� �mB"�>��u�׫D���iL����E}�T�t�Q�H�#���L���up���f��#��"Vtz�2C:3��o��S�j����Ed���Ckt�"�h��)�"՜�����XHNzk�#b����tt`������]vޗ.~1K�ʫ����m>M+�|�>GZ�=�)1�λ��g��\�t�c�I�3����F�K�ܨ�u������W�L�>��Iq}�B��Q
(N�����X���׮���Da��J�Q@Â�_dV�>���=rz`��*�4$� �naCҿ��8Кl�#���Y�#��RE��D�H�xd�!u��
Z�_���\��Bx��˻ �>:k�o�-�?����6{�G-]ۙ�ЋQ	=w��?����1��������B�l݈dp�9+n���v���� U��@���<�#=�P�o��;-ld�"�J�p@���>��P��B���}V;-��q���|����cwU4x��LrOHщ�Q����E�kXh|S��Ԇ��C��f�!�_�(���d���v1i����n'��)k�	��1i��U��-F;����,�{3�q-l��|ĭ|z��}ng�h�x��UW������Ce��Mӂ��fW�E�K� ��	٠��8��}��-�2C��2������Od��H��n>�m^�hl+��l���K��Z������l���W���>��,�d��!
�.��yÚ�А6�
"�X��1͟�p��YQ �"m�W����}-���4���m͝���