XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����
~u7q���߉K�|�S`�[��cO7�)RTf[M��"ʍ�bG�ͺ�����ġ�\q�J�??=��՝ܵ#��s��G���&���J~�قTC��2�ື���n��P!�g�2�oà�����w21������\8i���ñ����=خxSt�D�_BF�v,&g��,*wx~�rJ�P���z1粻T�q�, ���,���e5c{���u��{\�����Q����#u�67kήR�ʺl)�i��h �AxxlR/�U�y��]����V����QC��P��:U�4ϥ����y��[Ap��2q��w.ZhU��)n��QDK����=m�[Yr4�2����a�7��w�u���� B��u\l��N2�ŀD��{4���}x�eM�����w��6�w��qxU��Ν�u:�_�t6�zP���LL���v�� �q��8U�&�� ,�^��l�&���9d�����4"b��jgby����OV�)e���w�u?]k.��* �?%��h���J5��D�sQ�E1��
�zr̙��ƆoEBM�;�Y��hOa� �{s�N�Ft����,��{g�?�[/�?�ւ	��.��Vrh�#�iz��[�J��.�u�c.MY8��U�e���UOK�+�!��~��-�P��t�m������:x�;�5կ%N��mѢ��miu�;viL6��9���L,z\ �X����Z��^wq���a�����1�A��8�H?�����2XlxVHYEB    7265    1660܆_����+�}����U�N�P����|�b.��Hߓ��r�Y��bR� 4�Z0�!�0��FP1�YYK����_�ݶ��R>���3�^�?���`��3t�-�J�4��Z���y{�3���]�9�*��L?SG�`$}UE�� gB�w=с��e��wE-Ŧ	���E�}��v Z�kxR(����Y��41�$<V�d�8Cu�
ʔm������ѽ�w� X9\P0v�����,ӈR��R�	0�j?��y��.;��1�cl��OsI�Ky��%WZ�[��L��툪�T������v~��.�Ţ�����>�Ѻ(����b���Ə�	)�@C�}q\i��:�g(��~��U��u�"ҲH|���,n:����� \߁�+3��� <U�O�'is�Tb|4�c�t�Z�h��d�ŵ�`(o��,�+@�rA��Ն�ڋ̎A��7��Hf���D8���� 7�(^�J���Il��xӊǉ�F�
�z�
|ŕ
?�G/��֥ƀ��xxgv
�n#�鹹��eA�tV��.5/G�ZJ\Ν�Xc�����oŮ)�VC��l�{'��j�����' �t�ÿfK]	�4Z��욃o�s52A֙����{�	.�պ��[S_���������p۵��(k���D�89Ɯ�>y�,��:����j�@����w2%���Ú:�"s�Q�,e���0�G��� &�N'�a~����F�w�Q���[/�y���D��1 =�a65C\n�vgN�[ҡ�U{+�>�QI6tcQ-����)��p�5m6��y7V��)�볠�ƅ[N:5�0<l"2�X�D��+��N}H�o8��o��?vz�����|�������H����N�_ȒʫG�{��^%f�{o�f�����Y�fY��ʯ�E�G.�k���\���E9�8��]��^���U�*��@�Dh/b�A�(~|"�NDa�B/��ce�ֶ�!	�n��_�I��w)�)~��m�.h7-�t����<(g��]&��5�&�L��V�9����q[�کPKl��Ѷ��n�+ꓚ��G�v��1�:s�;.K���ϴ'�hy�`�ddE���G�|����/��h����t!#���?JN��2��6#�L�R�嬖�Х���Vn��=6XyF����-�l�+�xH�^�cx��a��ꮎjLAoAd���3{���'�}x�H|M�ǀ��6D1,0<+@���[2�t/��9��zj���:Tz�>�G�7���0%��F�����DH�\k,O}�f���C�u�IeV��u �p�H>Ga�ͬo��5�fB�5�`��Fm����D�4�����%�!�h�uPVOLܑ4��ڢ^�v���f��ە]ǫ���!vE���_,���b��q���Z��	�|�>YC��c@k�ty�ѣ�Q�	�㵹i��o��A���KW�n�V�2�A]�E���$��JO���w���s���T/�mD��v�N5��0�5�T��n�$�[��8��W��-%�(W�o{�~慻�����az��p����*�N���h4��0��
���;v����Ɉ�l焬G[Rp}V����T�u�d �
��Y�Wh7Y2G��G���=����o۫�`u��4K1]��n+PgRf*+��EG���bX�xp;�$��O�
�"����ß�O���((,�FtL8�,~dD�aC-N��s� �;�*H���*�����1E9/���a���w���?��Dd;�d�ޑ!B���������{��:S��w,z��(���{�}iF��'p���Ӊ�K�U\�`;�LT��B�Ih�ٸ%��-�Hw ��d/���ƀލ�Z.�:$pfbs���lR!1Q~��,8�<O�by�f�fVQ�lI=3�R���)�����P�4�)�����#�5X�~<;ʀ�Z�©N��/�_LrJ����%ki���v�6^S��f^�܋�b�k����;��)�&Z
��#�ߪN[�?��cA�fX�x��W��]e� �h��<Ye�Q��BGW�V�2>|���^��[l2��H�6�Զ�z��̍��}$��/WZ?�{����*԰�T��n^h����Ihq���Ir��ˇ %�t�Ğ�"}1ÎY��#!m�:�1�S�:̄��;z�OS#C�a� 9/�V�D�M�Ʈ����f$H�f}�FU�|�3DCA]������̝/\K�X&_\vS�Vg�c��}�+�}(d7�:yNl��ő�����?Jt���ޖ�M� ���8/H��/�1�spZr5]O�JJ-��U��;��ͱ[f��~M�B��;���B��d]
o���X^ɾ�$��5����S�M
"^�ݱ�Z�N)b���E�ٶϪ�ٽ�v齧`s-D/T��Υ��R1�y!�p.${^��`�ۼDRׄl]�[M�zX$x=ds7kG>�R��Wx~Y�o>ma���3�Ԫ�WB��n�	t���ǿm�c'#o�	ױ�X��4��A���	�Ps�u��|�L�Z�|�)b ��o��A�a�:ϻ'/�,�$�r�vZŽ$>#�F��%K�Xe�ǭ�@z�NUc�
�^m"��yy�"�8��JÓ�0PA> "6'Lk�pk�bcg��R@Cl�L�����v���#
�TsE)C�Vs~�m
,���=cCF���GQ�����klk���>���c%���4 ��#�r��u�vGd�x�E�E�X�:��i`�-_�Uo"}��8WL;9������D��6�S��+zV�x��W�t��9M���QN��ŀP�de�;U���2�`I:�r�@	��a��l�tp̃Q-��槴��r�=�dm�	��1V�L..e�K���L��u�����q��x*W�9��9�Df-�KV�X����`4�t#��r.���ài��c#(�e����q-ļ�w\joҳ��*D���q>!en��汷�FP*�cd�R�0h�Zղ�z���|ۃ5��9��� d��BX`��_�Q�k�*N��3a��������>�;!��y�K��cp���)>���%�Ҷ��PR�D0c����@ZGz-5,��W٣����T�`R$��ba� ��xeA�$�xs���x�Ӑ���� ���v+x|!�f%�v���>hl:g^��%wFx!#0�^f�깜�#�XkL�J����a��*s@N�I���#��|�g���� 88!t~�4�-+]�ࣰ!��r氜B-���k�Z�E���Q�J>��dd��&�/�
*p���Gߜ�,���6�'��
�%�;w,F�}���tX�-�T�����'��)��6k���9$</��]���ĈzɊJ?s<�X�7ɇ�M��+6�`�+E�7 �^6OM#����e�6���c�}fy!��/-՚鳤y�yg���k�_��=��Z,��A�������,�*�F����MT�� ����\�ŏ��Y[e!�Jb�ᔰ��nkcK۰���e�M5�1��#n�y��'I��9�1��T�yY�3��D������Fh�jL6
��H$��R�m&����3̡�)<����^1y�!�^�P��VF�QX9����bzb\�Ӱ��Ƞ"&�Ud;!�"
O͝���33xſ�cAx�tq�:�>�-yS=��t��%|!��b�-��"��G�p�͠;����5�����)����������=�*<6a�^� �uDGnoqR�T7�n\py��7��r|�e�*%�	U__��j��9��W��2x��K(z��~ O9P��dQ��z��@w|�"�&Qk݈�ު4m��N� ,���S���zU3�������[B�hz�������=s��Ya>�?��eU�ZI���`B�`=���ѱ諷AU��:��.�.H���s�Љ=�%�����8�c���,~D6���ݗ�[��֡���}OhP�Bm�T�_,��G���J�S�廅������$뇶|���`KI�[Ԫ�i��5$ܞ����F ��S����z��OM[u�H=��̘�����.l���|S^:��,��/pR2�G�;�~� N�r֝�Ob���K�wF'�rN�y��Uz��Dct:�_
G�PA~z,�L�Ӷ1iˤ��??�̗�����bO7�r7�қnP)v!3�a�I|����0�:�O��Y~Tm�z^�����b�ɱ_V���	)�2���h�QO���G��N����"͹Ruf9K7�k�Y�D�y��:m��%}u��^����*=���ak��Eե�ŉ���$��2��vh�§��Z>[��H�Ŷ<j���As�o�G���*��[�i�!�<0��Q�'�w
@Ѹ7���G���O��I�߁�� �e��K�q�Z�1���c��5���y�dR�[�m�������ON�ӢsgnQdE+������K𰲴��X�w� r��[�A�|O?����z�	u"�P����a<�-a��h	^;��Uq-XP����kܯ��I�Qe�����T� �{�E��H��%R��^dj�"�,5ݢ�ہ�e��B<���.g]�*��>�b3��Y��5�k�شH�٪�Ѫ���l���$#�m�.��V�l����x�ǉ���g�(�s{��,rAZ�`ޕ
�[EIn��~�J��x:7҉c7�P����>��7>��Y���k'8R�+'��^�H�9�Q$O�^i?�7�����M�����W?��O�1�(�b�[(ݓ�UCi �5�ڄ�pb��HwqX���β,ɐ4Vږ|�=슾�_�iy��_���ͅ�JS��UWh��0,++;�8L��>A~�a�]�h���GĔHO;�L,"�9,�V��dy����M����+F�<���n��	��!,{|8�R�=5�i��W0�����J��TZ�m���H��� f�e�1��z��$�_Zz�I�EW!0җH���R�H�[h�� ?�m0���7����b�;%j�o-:�jr˔(�h��_�R\�_���ޥ%YG�Ϻ����IP�թ�#*�������㐁��*����A����/~�:�_т8����Ӄ;�pr�j���Q�2A9͹nO��S��Yk:g�nh-I�
�JVn[~/�ۊ���>��(��{|>�}O�E�����Ip��b�'�o؉1r#�j<$w7��f	���񪒎_D���j��x(���JWu�_͞�E��Wt�HI���и�����(��%�XBᎱ �� ��b�JL�n҈E�pɱ�]3�Ώ�+��^�+���	�k����z�����+#;��rR+���$,�_%�@�S�x����$9Ώ_�	�[��eB6	���Ax�_��`N�����U	�Ԋäq܆.���隐�/�d�����{�V������m�����S�-���f*���U��_�(R��yJ�~��}��Z�o��I3@����ˀ
n��V�P��h���aՈa	&�pq�w��E�̷I1R�Y��~��<nٻ�Й��L`�џ;�=\�`�4op'��)]7ѻxP.4A=������a4���G��P���ݍ�����E�(��e��Rj�s���Q�G� �1��u��E��Um����fq$��-Êu�aymN�80���Oグ���3������D�+v�P��DN�gf