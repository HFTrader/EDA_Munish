XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���n��KjX3�R��o�2�Uq[m��� %��xk>s;*�y�e`�F�����̹�ש{���yrM�8�����}�<�~�V���o��YS�dv� �n��^���F�=w��t�uz-&W��<] z�w��u����C�PqGY�#�8�?0���:D�OX_Ȼ!�z!��r�-u�x��Ls\f:�}"p��Fpw��j�(�B�SC9L<ɰ�.�Da�� �%4�Ë���~��nZ��c�s�ם{�k���Yo���*�I���H���arLK=vwp��N�q� q���2_��q�Cş5�_.�&^K���!�ع�K�@(H������[!ɟ���'�	��=KSu�m�#�������XLtR���ME��њMy&���6�隀������� �ns*�Z�x��?��2,=Q���p��y��:�5�̀&����%�X|��n�Ǣ�����z1y���3�$���E^���9PA\_?o>NR.���A�[��������
�Rcq�x̀㔆~�j��Qެ�#��?e�3������ewB�O/�Q��t����������0!�ӊP�_~��aU�ڏ��U��O]{)vӂ+X���ʿHy��>�-9���f�wR^�!�wb�)��U���W�9413c�,�Q�BM�SV^��HvM����C~���(��>"���g�T��k�d9�Ax��:��дDB[�vh햗Va�|łayN��0��L� y����~���!�����T6�r�5�Z���Ӫ����XlxVHYEB    fa00    2030򷥿\1�x08��ڒ�q`�$.8�����:�~�ߖ<|��F�R=�&O��%��d�OgǇ�\j��!HŇ$)ğ���v�?��lNē�c-8˄��AU�:��:Nʙ�G�v�n�KZ&u�����{*os�'K�[f�Aiya�t�%�o�Vۃ�_����i�PT
cz��߽�1(���g@g��_:��9n�S\?Y��P���j���G�-7�х����W큦��Jז(��Ӂ���(�*��XcHn q����D��M�\��g�wa�P�l�J_����@�g����4�h9�?�pP�B�p�v.OG\���4Fk�!y�wJ(K,Ҕ�<$ٕ�^��.�*�̦Sk륡5��FV*���[��Ȕ�"!2>��h75n���*�5Q`�n�p��;���U�V��/	�Ӝ�>vr�|�F]�߁�ƉD��ᱎ�ܽ��P.�64^�6�/NƔC�| z�X�h��ig�b<`�Eh�K2����p��R��*yV"��$��2�s�=/����#��������=M"�F���(�:�K��Z��8$v�ł�Wh���~[$��i�\���B��� %&�����
d��ڔ����6��N�I�NM���+��@�
����w.i����^/���-�O�H��E\]]��� ���1��sd�lIg�J�mQ��v��uUAŸ�p����� B�������Z��SS�Z�+�q�+A�S�W��?p&F�p�MC�tX������MxA����a֒�Ux�iy�����r�5og�w-�!��2��9P*m���	�cۘbe��z�L�<�
�?�ԑ޶�A�:�bx�Vɓd��wT�40��z�'���v$�s�����vf�'�
�k��Y�6���7�q,eŎǅ��Z�X��pX�*�+r%%|L�)f�&�"���`!�P����\�Zk�.,b���ɼ������A�Lnv,⒅-��y�X�м��o�L觻.�3���7S����,�����B��*(2(Z2�A�O����p2��,o�}�Vb��'�xR)F��3=GCL�+�9��tZ%L���oߡ"�+W��h� ���j��R��0��J��-l�:�g��B�+�	�c*.q��d5����8�34܌j ��蝯g�q#�g�T�Sel��:R��(��֭�ذf�ý��wW��R:�dTV9#7�/��D�A����vrR�b�[:�m�O��j�x6l��9߆���z������o ���� +;�<���� $`�`آ0������ݜ���� ?*��ZK�+��*m���wv�뛁�k8n����b��U�ԗ�\�_\����]4���&O3�i$)-]:@��<U����HT�^�2V0���>�'Ν�,Z���r�n�A�:�?�톏��l�W�� �1J�f��)��RN�k|)���O��&���w��8U����=
�F:#���xr���ʝYW��Ϭ�R�k%)���.�L�.�X��-��\����Q<I���(OH��
�_�BƧ������G#�&��e�E1Yf��6��8YY�Y�-�W+�>o���}�&	r�&cw�QGZ��=�y�_S������{p��KP��6R�r������`���"�S�E4^��$K��l��?r��X�Dd�|���q��Z�?XP�c���i��-Q�"��jрt0��xz�@��X�l8�q��+֞��:�u�_���^2�IR܅3ϭ����wB�N�{���������}Ք�	�X��Ѷ�<�k�5��P��T�j�.:�K���*S[$��JG[�D��Ɉ|;Xd#o�	��:��������x�Z�*��xS'��A9��2�C*�H�v �b8�/��}�1�g�)���� 7�glm��n7/�NBO:	�fǞ��,:��Q-G��o�B��Z���An�V�Y̏ ���E#aX2��e�8���[C��.��)��4�OS�U�x��j���kQ��\����ˊgy�i{<~�	qX`-�3ه�4���
�\&���+ԝG���U�粛���7.+2]x�]x�����!�قQ�٪d�)�αO�����>,��e��V�R^�@��;W���$�R0b�M�{�=����f8��.ؠ���zɃ�b����{�������X�8�u���FT�\sx�EK�<�����P��q��R�^�	��>.&��3y���[1�`8d���0�6���,C
��f���nu]����Fi��߇����l0�Ǉ�'G))F��~����N=�'����,֓Q�	�>$L��j��$�&Y��2�
@�T����xDQ�SE�2Հ�K5��t�/�_���䇇�9W��6eI�A����B�����=��)��e�<G�������5�$�������������n}VJ�+nY77��%+��6�6�/��nIQN���&�&sz2�j�OR��u��[?��;;[�at黕p���7[��k'k"m 3m��5�*� A�k���ol8Z�������6� R0���FԌ|9��x����$/�����(t�!|`(�1��t��[B&���]6J���y�j>Aҭ3�@׍�31L�!�� �c�/��J?OC��z�$���M������ߘ��o��b1M���2��+k�ĒӳEq�H���͂���[ǃ�e(���|6�L�eլ�q���C�Y��^�Ƈ�Cj��8v��}�yb�s����6x&f>]�]<�D�� �Z� xz�ں
G*f�'�B�hs�ț7;�O�d E�N@�� :�U^��y���u����ut�-Y��\ (4�i L�r��n؜���~�αr#4�V�УJ&}� /�1��eG�me�s�g(R^�U:�Jz�T�!��(�CpLS����m�[xضb�N$�؛FM�X��pfO6��E��*�|����3��'��:_~�h�5��!C��g�%���n�[�:�����$�v|,�ꏄ���47*���lL��`c�k���5��c
o&�/��9;&�#-��I�dݫ�u8&�g����iD�n���)6(��Q\E4��j\�[$�Q�Os	�ɍ]��=����w��n�����9ܯ�+�r:E�_I�(�E��o�z��ި��E�]Q������H3[����؂G A�t�?%��fH�?��w3+Ȋ���Bu���d�9�e���|��iF�z��`D��SG��{��n�,@��H�dh�����c��*7h$u���qx��t�%'�u��h�T2�a��"/�f�9@yY�y�%�w��ݕuHK߭7�t��7�q�M�ҩ��\n{���0-ՌJr'���b|�͐`�v�o�@O/�8�U�x�w�-wy�As����m�%�0���}�;`�IؤQ�j�l��o��P:;[�b�"�����.��}a�JZA��>�Lij�2&�h�4t�܇�2AC��ۦ�pU������Ћ��7��AVs%�&��>���n���rT��Ky�ɓ�~�O��$6��`�gpm�3RqI��b>׼�٨��`Ed�g癃#œ�[��]���w	^���e��	+��z�ȩ�1C�=꥖���*�+�n�B�!���v�s$���� Ԏ��|�m��2*;q���|��j��gҦD���4{���b�g�ow�'��l�z�7����4h:�GxX ���:^����c����< ����\�H]�u�@�8����{{�|�L�W�7�xY��+>��r�V}ek��K��ctO�n�;�������;�C �xd�5@M����s3�JU���%���?&��=����;�9��R���y5n�q��2� u6ŕqY��Q5����E|�i� ��Ϟ�.��P}TOI1(�����A�/�_�:�f�d�AB��Cqm�"A��Bu �-u�|�ዊ������Mn�sabp,bq�&�� dЦ��N�_�=/�=i9�L�gXeġ+�c&�v��j�y9��F?>#�ee%]B���J�Ճ���v�qf"�;�(�\1��zA��k�U�ȱRs��Y/@ܻ��<d�=ȼ��,�o �O� �1�l>�Z��l��=�y�ύV��~���q9���N"��
��{�M-���iz�[�z|��߁v7��ӵ�7�KYӋ���]��rw=�K\�x.3+��)h�l�d�$Tv�Z���x�|,�t��F��^��a��އ��ߊg��ˁ��FK����!�@P�?�V�f!�kx����w���>O�*I��_q�9�{7�
S/; �l�0Tz�y*�O`��a-]1k�|N0�;�����r���Jt���RlI�!�ҏ�ܱ�s�?��ZNT�4��ԑ�F�Uj2��>�F�B�ֶL Η^� R����%��*N�+έ��a^1��0���QňܓCa�p�4 �R��L}��ADq ���U�xv�F��M4��k��Kc�W�� G;�֙�K�=����X�����=f1�x��ќ7���	�@؛=�����_2u����Ed ݃o����l�v8~�*�'���2�$����`����$�4�g��z	���ڒ��/K�}�i�'�)U�,�&�6tދ�;u�_[G$��X�}�P W�L�(L�
�z��pZ�>V��Bņ��`��ǖ[h��%�a���w<��� �%�\���qj ��~�s��DB%dm���#S]^Kgm����� �G8�l?�|��fف�+$p�o�#m��ڊ�A-����'?g�"D�����͋��]u���ߤ���I��򇤇H i�+��?�<����Hb�6��}�d ���_@����Ϝ-
����4����P�KF/pY+]ַ��O��1�ں���w��$�F�vL(�Ζҏ= C��'����SCZ��x�im�4杋:O�Z<�:�3Ҩk���Y�K�(j�f()'��of�����'�d���B��3 9��0m���� �����Х��~��%z��u���:e��@�";��ɑ�(1�-�+ ��!5�{����e��/ޯ3M�@I�t�KD��N.~(�(m�ZD�n���Hy�ݗŅރ�p�<�)O�[��-���X��g�=�t���P!�ݮjÚ����1@�k�+e�6�L�1���K�L���p��nkvFT�V�9� -��QUݑ: �������fG����8}Χ~�Hy�������zC�mL,�.��4U	S�R�W u�K�77�j4�3uy
��z�<�/��Y���;�z:~6+���>�!)���� r���H�g���hF�iT9vt����U�ĨJ����O����ڭ��Db1e�u�w���1U��a�Ͼ������GLsƈ��dP�^��V��5�#�߷;u�:���&�+<�-S�*� L:����l�~�Z+�]����N�!;���.;�r1�Ӈt����NK�����1����or.�5#�4��\������海{�����>�1Ub�x�|�! 
���WdG��m�Xp8G�Q	)9���U��-���6Vy-�^�}��Eu�{�p�2.sz�D�6cL�&��7dS�Nʳe�]��׍�� T��UF�����*�u5|K��_|��mM5�1`U/�Q:6*�3=Y{ e�Q6myi�]�I=0�s�w�A4	���������ڔ�i-�H�h7�R��`�X�8�Iǥ�6�4�E��*�˩��U���������9$AV q&����+��Nv�z���
q�l����4{}2�8sn�c�TX�,��f��J?�A&��c����d1�X��S����5�<dN�y��
�,R���	<��+��+$��@ݵ3��$2����n����-��Y���I�P^S�rk�i��k�./��ޗ.;�4����t�;��������v!���rY�����~u0��kKP#�)ʂ��OC�U��e'��?��vG
+���>�3�ӥd|t�8��%�C9�yl�|�sy�k`�\�Z.�0��Y�������Q`����Ѧ��+��ñ�0�"�H��-���*b
߆��L�#}�i�-���/�����M	D�p�����Z�#��ʺ��sS�i�w�wׇ��my�#݆4);Q�_�[���C��#h/���(���e��c�~��t��ݖd]0�@W�Ӭ\9�S>ރ���6F�H]��i\`�W/d<�	Y�Fn-}��Z��G���E@-')�L&�;�3������N����b�$��'zO2^6x����#�1��X{�G:�N,%'��#S�<�G"�p�V��xϧ߀t>]J/;`�v���e(�0v9���8]G�2d���:�kM�*3_��B��*�fJr�`4h o�ep�k�4؂5��	�:�4�O�v�:�?�1*(9���r|g�g�G���%��ԅkʒ�{ D �������K"�n�Ik�Ȳ�}���l��V_�{���|���
c�tu�������ڶ �Q.T��&!���U�&"r@Xq�~�Vc"�[��6NB\�3�,@���nZ�Tdw�C���w'��9��
�<�W���Ѹ'?�o�ï�d!��l�-c�i{��y' �q��7W*B4�J��:����T�qo�QU������*{�%���3%+�ʄAu������!o�� ��߀,�bf��Xmc�*���}ۑ����4��1'oo�����$J��@��>qR�q7��n�Y��-b�?��)����G�C`��oK>
��~@����� �d��ƀ�\
�]�4x�yK^�n]���e����u��/�Pj�����B�0���t������Y����:�V��[p�rm����0��@�ځ����-�H�Ӝ��H�VH�Z%�c.Z+��h�R�=��k�	\l�(I&����nv�%w6���'�u) ���q�l�b�Ҝ�`�����~�$���iO������FZ�Kp��z�QQ�wI��qXb���<ǳ���z�j���Ca�sȆ�Yᐠ.�-��
�������ҹg���͏�O��q����m�F�I��tZ��ǉ��*�< ��r7�Z�j��3<s�NrW�˞�x�>�F��A�N�	퇝����wEk�����l���(_8A_�ϧ�I�[{������FS��Y�����$�,�t'�w��%���(�ݠ�����;@�̕
`7X�� ���V��������Ⴐ$.]A`�k�3���`�o!��Hr�0��a���ʋ�07�`������ƅ�+@N>�"):
�Q&����if�S@��uIK�BXks~���+P"�|#ԜK�0
JBg���A���X��*���.Y�;����iP0�=�S]���[�a~'���򲓡��s`*wTy�@t��.�!���nj���G.#��B7>�4I`n�s�^_��٨�n���dIZ͝u����, .M�+�>徏tϴ���[Ҹ
�cgi b��C�l��KxI@���}fv�'�:~���q�.q<���E��Ϸ�s.�g�d���c9��B�6m�>�J�&9�~������.���F����Y=�,����N���^:V��GQ���"?J'K#�k�;޸��P˝�kZ��M�ӄ�q)*(�)�0�hq��;�j��GK� �e��b#B{��X5!�~i���²���4�����")��AWQ��l�?D<��u%�H>zi�ˬ�!8���c�+R�g��5���U�u'5��>�T�i�%x�0둵��Oy���Qi��=Ε{�x���h
��^C�VE����n'W���d��O��zG'~�
���k���m����߰�5~B��{H���v���*�kl]5P��d�`BL,o�y#P*
�����EF`\��Y �mݾ$��]�o�Jk��
�K�$��g�8n7J�����={�/\ZV�N�V��u�e�ybZ����g��Ғ��fQm��'<@^p���D�\p��\��V���R-�F���w�]S`�r� E�S�\/ N�Luo
�Z�GD�7��V4��@$�Jt�H@�˔���_5j�20��1�8ꎹ�v���}.�� �[�Bin�Z�%ai�5�L�����_D������"2�d	��n��LN�D.�(��Rxb�NXlxVHYEB    9620     d70����j���s�|����ܨ�J�$�%:��-��V�a�>�N�p��P�V��.(�z�
s�7U�q���"I�K� ��ЂP�[/vJ�wϬ���˩�����Ct�-He;j��ܧ� +�r=�>���&��� q�|*İ7��V���B�|"�Leo���c1ks&��2+��e��� `QJӿ�Fq';R��E"���W����s(��>�:n��Hj���%R���;=r %��
�ПÉS;��$��	C�=W�ۈ �f� )�x��o�R�c�)��5�� Ӆ_Ʋ������p-��J���H���� ��V�w���2F��_2�H}L��6�Tf�0�����6�}u�0�����e��v5:��?8����:M�yrU�4�k���'�gZ=����"�˛�G�{+S�{�F�sͿ�(Ϯ*��ԋ-��$��YcIJ����%��-f�ֵ��c�V��c��=ّ SG��Qp2M��GO9;�%2��D3�s��,k`@!�ϒ�zr!�&t r��+.1�K��Q�LAt���%���5�ϲ����O9~�55,�s�`z�
�ϡ}�-�t1�FV�k�!�*n-)c��ӆ!�뇆���!��>��z��:��3q�c�HU�հ�7f̄Ĳٕ��2���Q>�U�q���J�A�i���^�s�{=�2�,����8����,I�h4H���o�5Z5��v�/;�7D!���{����P� �mkG�b����Zw�B�� �k8.W̵�t��Wә�'5��dl���x
2l�,m:�jK�ӂ!�ڇ�a���_|2�LM��/Ew�����x\�CV��LD>zNV�k��3����y4O�����Ɛ�BQ��Yx�	&9�r=��F�3���b}�x-�+(��,9Zs�x���g��x4����,�|1��{��5ުГ�r=PjN��s���R����fb���B��m_��l�L�z���.0¥����V��.E���~mhY���"<5ޤ6�WU5!$�2:��@���d����p4�<$��e��/&���?�K�����R2�u��|��QP� vQ�b���^ \���Eߜkb����A
���bW[�j��:�����<q��n����ֶ��K���:�xL��v��v�Ȩ�"v՗���<_f�Qh����m����c<���C�VPJ�x�1U�u%���0�m�E�r��5���8<��܎��mԍ��V��o:�AH;�#C�w�q�ZXkN����F�ě���ߗ3 �R����u���L%H�����`�O������V��Η]�ݹ�as�^߁L]�]�JߑS���X��/7�j��M�;��ZT[�f��_���4˵={Hl0����[�`6�/vN�c��;�b��[�g:AJ�t��A�TL���E��X�$	k^���1�n4�*�p;,��)ZvG�ä�zq����¶nl�/WW�c�J�;��%u!���휏�:���l�8}��T��ty������^�Rf�]�ӕС���DK_~C�}CNO7�[7���X/VWZ_�u�f�X����-8�����x���n@+I͢�٤� ~|���mڏ|��.����_��E�m@�����'��AG�N��cu�>Vzg�mV� x���tw�Q���/Ho�RK%�t�|S�c`E��q�c����ro�/�ϕY�R�%�ޱt��B�*�E��} [	�qIe�W�j��#SJv��N:
/��J%������/#� T�6앒dLh�5��8�i2Y}��.���tx˃��N�$@�N=�jX�r[��b���1���(�b���
�	�3�2;��k��Q�u�0�T끯�MW�lC������ ��=��r�ޏl���[%�wzvN�����;qh�U_��_��c�sM����~�gc�g��$C98d-řH;e qS�$��L?ai���A���h�dU�(��4���`Yܸ �H�M@�a�'�|�K<O��!�Ix8U�-��e��X��8���Lu��`���%c�3�4��KP?g��WN.v�s̈zҡ0�'T�N!����T=���C�}�t���.��r_�����i����}:$�d^�`Y#�����ŭM� OC�?�AT"���21��Qi(�&�z���x�>G��X�aT�T�i��]x�]�q�.��6K�[���� �v�I;d�Xϳ��^�[�΍�X���04�,�*F/7�y�S�e���xa��#$Í;v���舖����??�.��x��f�ޠ�Hh�{E��hV�J�fr�K�����}P�.����Fp�;<��5��GW��&�B�������7��Q��m��UHUe]��'v_���ʛg��
�Y��"^=��Am�}~�%��g���eK�x޵!�����P"j���e�$]���__�C�@k(u�F"l���QN�l�i��e��̮��m!�9�SH�("���u\��O�/��*%����U�@Ǆ(W�(I�|�W[��VD�Ë ��i����o!���8oZ�V��$�X���� N��-{��nOދ��Q���N^Q�P�Ċ#0�^�/J���zp��]�ڼ�Gq���be��C��R�/o��h�M{��<�Z���0kL� �;��8�����̏dUˉXX	F�mF���L9�����T��΄{�1��Q�t�s�Vk�,�l����e|쾘ب҃�/K�\2��a�Õ�[������vy��-�&�!�Dzm�z����%8Q�T�{��"�k���2��<����J��˹OQ���(�����-��³�'�:jyC��*O��˺+�#M��0O�١��s�h��5��.�>˿]|�"h�/6��(ga@Y�"2�����$�Q��j��S��J�ϭ$��v�cJ��YRn�2���ϥ+v���c��w�>�{Kq�u�����E�3�(��x�3زaQ�,!^�_$�N�6z0
Kj�w�<��}5�\(�h��I�yl^L���6_����0+�p ���4#D�0 4�)Ng����EZ��=�~��˘�}? EK/�V���to�o���{�=]������� 87��@p&��~s�J��+|���`M]��;�>���tf3���>mN^��7�k̀��r�����z����ֹ�rb�U2���xT�Ů����8(�`�ǻU�Q�<:���8�Y�4���á@>� ���d}鿮�Gt���mS'�5���.��@�D_���q�P4 �,x��0=���_�$��7���y�	z�SA"����cH���e�
#��.=3r��
q�BSV��M�慞(R�����Y�)��e(b[�ͥ����4H۳��B�UB]���f3�H/y�u5�������