XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w)����)4���e5aTU�%Y_��`�}���+�9ǣ@q���)��1Bd�j�0��u3��6ĸ�aX��ӱK����iP8蝲&�Z0F�~^�B����3䪖��ۋ��^��;���~�ߞ��i�uю� %-�K#Fz�~�֦7���?_V|W�Dv�����Tttt�L�_{��,6����\���C�/�X�#��4�U�뭖��l�q�p�=V�Yʉ����Ler��k��&�P0u��0F���!���Ȁ�;��yu�-z(^QK<�X��k���hU�p�xN(��~��t5�������rnK"�7���lf�|�L��r`R�fK5_��MV���2�v�8z�\Aǥ׸ZG�����x��	�{��Rr�y���A?7���\��n.�
�{#{�Z���T�!y����p$4<�xR�XX���_�Y�.X���iн-��Ovm�6V�n�������Q6�C8��GR�޽^h&i��c%(�Ž��$�M��;�� fq:MX�~cʞ^,��,�[aUyH��/�lA�s��^<�%#�&,?A��q���	��Qviu�cW�+W^�('KTS���!P$�N�u��-㕮���r��7Ac��H�A�eYۏ���!BdG+��4 ����)��,��CK�-�-[����W#���@|<�!�F�n�A��z��-�B�1�~����H,l8�@�����Ŭt��LJyGl�.�[8��6�;|1j�{6�[��®9�V�XlxVHYEB    ea93    1880���l�*���9W�1
K��a#7X�O1��c=�R��`����Gwi��w4�u&|�f��i �#-�*�J����PۨWH�L
RK�3,��>d0F�*ؘ9Y	#с���n<^�ɬ^YJ�wH\ o��N�BF�Fv𦵙��y���d��r_l�Ȕ�O��@� ?��es���`e�g������ƥ�5����?�l��ԫ�k�G��6���U���/I_.���pd��O9��\0S��_����#'�{P��|�T��ҿ�}U�㲚+�������Z�ˢ9^!3��9-$Pզ[��U����/ufo�`_M�MH�W��u(#�}Q�c���b�qQ�WY��BsΠOCT�� z8�m��ot�e;%8��	���~)�75/��� S���@��t�ٖ�'� n���-�#�v���߈���5��|p�.��m��ʝE�����M�M( �ZH���}��Z�۫y��֕�j^��.����90g;���CՏ�����y�Y�:�}JE�/��jM������s�x�>X��n-�A�Lu��F��{��"�/�~Ⲝ��А��VM�<5���vxd�`9�r�ŕK�I���ԉ��hc�=�$�����>c�w�W$Wsa���z�!}JDSa\^?\mTn�*%C��p��;�~��"J��H
��*�P|h���!j��zu6<���V��§��2��|�{�_!���*|#��]��U�#��& �g�}��yY:��2j�C�=��}��2�A�� �_�����Q�M�X^��bk�#�wJ*��`�Ƿ�PJj�K�QQ����G2�d�����\�:���H	�<�a69X�"���4�g'�&�:�sx�+(��}>�����CR^���8�@�R�G�M�����P0�2���ro��?��;�A���4%BJ����3��րT���'f���a5�ԥ�q��f�����!�G�x����G�K��T��BiZ~�b�"�#8�d�a���jQ���#=&��Ҿh�M<1"����\L�v�U��2< ���)�Y�}}�R�|Lඡgf��t�x�r�䓶�YN޽����	��o?f<).�)�k�ͨ�:Q�`̧��P�Sh������O��B�4nqԍ�H��~�{����	9�qSu�k��h$3��NB����H��W�u�y�?6��Xz:��w>�MmSҚ͞��|�[[l�,� ��y�n���n�#�����3���@���K�õ�C�B�5qj��o���<���DtU)��bBB�?�`����@a��@U�-<n�iLl��I%n�]0fcH�P-����n�By�'�T\@'Ƣ���$ܼ?	���MJ,v-�J|�>�3u��E��m��5ĨO7�7�~�ٖw`͜��>j��l>HϗS�� a�cy���Ư���`�J�������o����;�3m*��!�{�VM��?����{�U��C�D.��%̚R��:a ��(X�[�1��!���گ�rm~/&�e�0�?f�N��`�H���$n�Pael���\�Ti�qM�v3�V�R�5k#�C[{�� 6����$s���!���N��胎x����Y�YL�]ь�Ʊ|��)[@c׿��I�}�瓌'��1E�2��m�?ѥ
)��K/u%4�t[�\E�E@1It��k?�V	by�P"��`�7L>�J,*�V�,v͝�x�[>;j���-s|lb4�iޡ��}�\z���8��?#�/���2�G��O���� �X�~m�Z��h}��o��u�W��4f��XXkeQE
Gb������1z�M�	�
4&���2y����i�y;�}��M����
,������/����v���?��Y�uz
�;��\�]��U��U��j���1��Xe�ُ�*pl���hL���,�g��J*jK&Q������F$�:�,6��)�z��d<���ͅq����42�w�ޏ�&�ܚa5�:N��9t�x|
b���i�&İ��[c�!.��.�ڽ�ᗮbPM����;�G�U��6B�M]�X�x�1� 9����9��Ǿ{�}X�왪&�O��Ⱬ>Y�(�>���C͌\6Ly(xR�}��������J��b��R�n_u@}{�*�@����k{,�b� T�4�Z?�hH���.�oǎg@��(����M�4]b�6!�
�TDg��#'���"st�򹞛vi���4b�v���(�Im�	 ��]O�J���Y��e)�}Ln`���9���o��b�T�gØS��ӷ���a-���ݿ��)o�B�� |NK�⮒�� g�������a��'1��wC��{E$D �H�;n��Fc�Buf�� ��m�ꓛ��2>ꎲ���N)�f�i{��a��;g�#����/ �᧴$��r,�n_�Uog���I3X^�9V�QZ���EN�_��'Ź N��{���\�A���-4Z�Q�ip&W\�[���G�I�>㻮nO~�a��$�h#��ɆxV]J��%K�_�v�
oφ	�qf��m-���=x&-�6�k��t
���y� 9� ��G�&`5i��u�t(�93�G�jlu���/"e�q?�}&C���b\�*/S�uCn��4��j�n�F���^�n���+.Z>Ѳ���W[bJa��<���=)�(H��YrS��7�CO*z a�A��#Ȅ���.\���u���,��T�������/�t���gP�H��Fr5��_��x<g�^����1��z�r����bS� }��s�k�,1p@5a��>��Ͷ5ɘ?!̅Ш���ER��{�AY�j�s�^{�ڬ��v������)���b&�|�ƼHL���{��_j�������Z�M ��?o?�`p�SgT��x�~'�|��3�H
%PX
8���?:Vj	j�2|�U�=�Й5,�*X�������b[&�^�1A�$K�M��xXEe���~��[ۿ��t4��~Bk���V���d\�-;�R��\�;�����P��*3 ��6���M��m��6�����y�=;���mX�\Im��c2�^�	p���<�M4��n\X���|����j�Ba�n1��wn�3�S�!X+~oL�SNO���_���o��^��A�&�a^����#�6=���ԍo��r|�1�؀e*���0��9b��H🳤�����2� ��s�_��Z>�|)^T���W� �.-J&����Odm H[1ۺ�ԕפǇ�.��Py�c����^�{���ɀ�w3f���gѪ��2��K̬I�z�Go!6A�xx�\��:T���Njg~dz�>&ު�H�y植��B���it3�q��0
CU��<d�h�Y�V���=PB)�wAsg����P�`�m
�Hf�a9M:�@�
[��g
u7�'(�ׄ��-y�aa�r�u�T�d�0&Իߊ�,w�!m'��i�Lk��&yS�׳7����H͢"�8B��`ݾ��U��s�JJ�"�9�͘]yՆ�[b�,�2��{90$|�J��L��|���]��?���!:�yu���>�y6�Ss�R|��ϟ`�[�}_ORo��9�t(�{ٓOM��}Ϯ�'��Zd_�u�W�$��ф�Z?�r6�9�y.��E�Q�T?�g��$�u�Q#�d��T��mP7 �7�l�l� $��.���d��d�"��O����xC���R�)d?�K�5q�L��w�w�{+A�q����"��H��5����&fؼ��5,�BH�6D���5�Ө1����E�Bmے��))!�#⯗��}�#$'j~��8�L��'x���շ�iS���M��RS/2����vnW0��a׽Yk��gw��o�h[F�xt�[R&�9YE{��ݳ���b� �/���M�2�>zb6b.��g;&��!��j��dJ�U��be�Ѵ�D�%;gB����<���Dlq�&�_}2��R\�a�R�t�C�����λ����`P�c����-_���
Z����
�+\�f�&֠_H�0Px ����w
�;	Ƕ*i��I��,oB%���S\��p���n��B}�23���'���߲^q;�h�ĵDH��Z�@�hR�j8�Sz[�Z@�B�3Fqq���X���V�@qM��03���\��N�E�$�e�z�6"��XLe�'�v�����[�-ER�c���_K�
EAL���O��dh���+�9�p}⺙�G)���isi3𴆷=r�)�����ۤ�+�ȗc�q�TPwV��1{=r�v#���_�ԋ��pJK�7?Exjar ��a�- �:�\e���rF+-J�j�x���S˜м"��x79+�#3�m:��V6T�)wR�c\��}0%���"��˶ȓ��*�u��{*&�7�lF�^����T���o\h�X3�*HHe�go�U�y*�����&-���x��$��Fɤ�*�)��㹩�D����*!��l�k���6�R�'�L�#�ٶU��pf|�1�EmQ��^2���}��߾��*��&>��c�*����%/�n���.Ii2]�1 ������2\x����I��:C�͠� ߛu\�JL���Z�U���P�z�|.j�G�+��k�2�4V�J���gt��ػ�R�J�����A#��r��8hfY��#��@"q��G%�%�����*����]�i�i�YbW�%�ii.��|S���~,p�#pɎ,) ������^p�#g�2�f���aI�ru���q6�6��v A@S)2��Q�g:86���3��fШ�2A�r��| R5Y)����=��x�fH�P}��%%�a�K8�o�̻b������(�A~4gj@R�[��v�F��VNJ����n� ��X:�ƼQ�\I�7�v%$��1�WǪ�m�O���4R��HBs����b���������uη��3���%;���M(B��$� .hsYWF9a6@P�7�IX���J !F-aL�,
�XL��tN�5��h����2nq��F�bR�����%�Sûz>�1��,-lU ��/�.S����Z��r
<?�MXn��m���A٦�U�i@f��m�-
:n�������o���T��T��,�%y[�ǜ�R�����ǡgZ��a���&#���!���e�UoOS&�>�Hb�Ҧ�	�C�]��������r�VwB�Z�Jpj&vݸ1�b��5�C�ث!�q�:�04��������ё��~�/��Z��+�~ɕ���zV���s�ǵ���g��a�h����%��h1�ٿh���/$��Qap�&�5`��i������y1H�c�v�/<��B-a��k_��<3�ê��oI��'&hr�>�x��%s�k�{[U����i3�vR�6�g�(Źd�"q�`t�jd0M��ֽ�J�p��z��� �R�.���C+�O ���wxQ�h��&22ɫ�"��TGz�h��C � @Y~�X�E{
EX��YSO���l�G�iށ�����0pۖ�TDgfs���ѵ�0��������R��0��?�Uh0�	�$��3$v�"�im���Ԗ`�!D2溉;��[��sk������e��#�1R��4:;`.`����*�e��c�j�,=}GE�(fO�R�_�i7!=*O����c���3��zr?쾍��P1.���G���<SMP��Ӏ��o��A���sKf��s�a{8V=���#Ft���6��Q�0��ʣٯ �yrF1s���)m�+:O���&�+¢�M����:孯��A��Wي�t��6�j{�Lu|�r�ʮǚ�S#���~C�Kv��׸"��A��ө�O��ԥHB�4�s�7�
~�*�i[��G9�
;H�|q:P<������eYb�j��2G|�T<�U#s����2�c��ag���X����+f��x�r��	7�u}yH����xY|�����7�����:�b�"<��J�
�?��`$8����{lq'��5G|uI=�+-�P�s�=���mq+�đ�ݳ���Ѕ9�c�w���Q#ӹ�Ý�5/xulj�(-�"���ֽ�l^]�W���z�{�o2#�竸@F0�r��m�1wL��7,�q��d��(��ΰ׶亍���29*!}X��=?���|D�aS��]�g��.�]���	��(zu:��$`