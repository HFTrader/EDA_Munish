XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���̐/�ʏ�/N=�ѝ��`�"� �6V���v1�b w�w���
l$�d�ք_?�ԫ�Q<B�h.VC��T�uJ�g�2���B4W���+rs�k=d`N�юl�� f�l��)�����/D� �f]D��WݩXđ#L[7;���D����/��W���6�Dw�D?�t{Ќ=�F-�n��o�|�X�ܟb(�c��
�ξ65Z�����7��������)�\g،�;��G�1����ߤPxhm���CB,y�vksSL�q�����	�P�"��@K��������f�'�Q9��e��\�����Ҝy���tR:V$��Pa�D|΁F;����&��m�ҟ~H*\aR\-�E[���LЉ�rp�0Ҁ� ښRe;ď�ˆN��_@v��Cώ��o���!�o��E}�� �9�K�h����:*�熮�y�//|�ޘE*�B"�Z�Y��G�Ԃ�(R��E�tL�T��ռN7��O�p�'P���*bJ���K3��3�β�5�4�YP�#��C/B����@(RL�C�f�މl��S)��sҥ���	��h	��d�I���>���m��s�F8���u���cL���F��JK}��u��iّa�j�9�\X�{�#,BA�����C=+���nҏJ��/!Ju�-�����+A��������X{�1�\l��F����������f��ِ��y�,)C�vʢ��X�7AO0n�@X��gD��p�Y�x܇;��t_Uw�XlxVHYEB    4a7d    1090̈"�A�X\�~���V�$S��7XI@n��@��a�M1)�a�
7�C8WJjR�&��1�"����ˍAj/:W������MJ�2d��	�5>�Ts�a61�|����F�9�u�;�S(]�\�d�;i=�>kA��n����Y���|9ή&�c�)$5o��.��V�l���>�.�ȧ�Q��*O�7�ל��2Xk5x�d�z�S��ż��9�{�)T��޸�R���(�#��-��D<P�
����`�|��.��?5g*7����������4i��XB*�?^�exx�����>ƚbD��>$��5���d���K��M��5��'yi��{�?&!aRE>uǤF���x�������lZ:�8�9'(w ��xS:S"�n�V��W�K,���;�WN^r���8�0U,�-��(.�UD9�K���"5�c��ҳzZ���rȇ��3��%9 �~���ka i���|��35bad�6�����2w�G�窞�(���Z�A
�&1�
=�ً�g�7�J�=��J�S$AGe`17��{��NT�B��d��zA�~ v�דv싴pkS�L�E�x1���.��}�Uf]$ �pq�L�����c+���U�Sn��tZ�ar �'~����F���~Mt$�k7 �/��\4w��c���x��UЬ���b�����&d��`R��C�\"J�j�d��Wd�0�B�@YV����� K��_��0{����Ī��<��z�[�4��cieG)�9qv�Y�:��4q�䃇����Ͻ�ح�4��4+�܀��NC}���}�[����C9�jy�{���¢_�	�nCquY�������CHU��o�Ç���;����"@g��	NJ��z0>��z���r!�$B�R2B�1>1���*���p릫�4_��-���t�'`�mS��zN�׿�>�p3�&!:��Y �H۸G��TWMa3������o�.8��?/�\E)�.�y>�I��3
���۵��E6�9Sx	�V(��<�����u�m��/5�k4�C���2�q;��ٗ��4a�����I�p7B��a&d�����3��_��R�f���h0�_R�|
r��f�S/�_�W�t߆�E��X"p�{#��	�FFy���<�s�=�T�ָ-W|}��~͊ܥ���jH5AId9֦�;<��!�Y0�}�l��5�f	Z�խb&�wC밷`�wE��o�=�?�]�"����W���2Ópۡ�8��5F��Tg�^����BjUo8%�A֓��zR*���&���eJt�	�p��~�NrW��(�]|�ti<hj}��������v�*/�n���$�/LD�+i�)'�/��cf�����Nvm(UHH0`����wDZ;�AzKe� �Ӊ�����$���$-��p%R1�z�P��.��Wz��=[�O4�!_��S���nR��̜�*��50�W� %%%��b��X�ۏ!&����/�F��)W8WD1��d�S�ۄG�Y�8d&����1A^�܊�(ok�6=�p��M$��8�P�^�-X[��Ӱ���o���"��=QZ:u:�� �X�G���&r�W������d�k�]-ĺF��:�@���i�8���TQ�8�7�Qũ� 	H�;�K��ת�Fd7$�$C;)�vf�Nф��MC�L��q��e���C����g'��T B�Oϔ���uV���I
5�V��G"B��?g�P<	$�^yw����@&�� �񋐞fQA�O'��:�_�v�`F�G��c͘r�$��j�RP�ա(M���ި����*2G+Quߤ=�):�$�$�F���N��G�4,�>C�2!n?9I��k}:ӮD���2�a�#�T���oj"��E���>��`��/�VM������}�m���K��eg�z�{ �!�8��2͟��C�9i�UM�z�}���mPϲ`ԯ�6���ؠ��F�^?'Ŝ%� 1�}fq���$>(a�0d�����<s�^�ߓ{�D�4��H9O\�r�Z(����4[�&Ub*��&�������J�a�Վ�!nt�ؼS\��,����2x�������u W�.��A����8e�W�=�����֡��#��K;oҐ�����0Ľ^�&>�������(��zfU�p���aB��eo�����M��B&ݾ��\
�E�w����JFв���!"�Kx�N@^�M!?�P?ږ����9Fdͽ�8����+~�ic��m�	�l�qW�9�$,��� g��	�kgSD�ͣ���r�*+�561+?�2���ׄ���v
�'ؘC��E�Jy�����1��m��!�mh�M؇�B�p}Í�) ��nJ��Ȳ`KLY�B"p�u���z�%�D�v�>KI�шr� �rj�D�/sloƿ���f��ӥ�T�G��ʸ����$x˥n����c�������jE�~/?��uB�)+���vJK�EjtHF���~�<�))Ͱ8g7q��S��ymz�2G��
a���-��Kh9 ]]̺�v�F�R���-����8��pHD�Z�kX��4=	�m���}Ԉ0�������|z00 �L5�_r95;�6U/U�M:�����&f�M��N�],(�&�Q@@��h�����U@V��(ђE�,���)����X��o� ��X��X[\,��y�Q��� $�t��G70�/Y�?�z�Ǉ���M<�h�a�PС�П��x ��-�k���'�M:O��͐��� &ɍI(䶏sޘΒh����)ؓ�A��I-6be��� B�1(���!�a	�M0D�h�^7x�����"٥�������"�n�w�Z����W��4%3��D�A�r��F}t�>��Ƒ��֧�1�+�@b;\�Z���4M�ח���,���_��;����u�z%�*LfX�A~�r�bL/�d��-H�2�g0&�Ь���w����Z��[��Mu5ߍ|�iД�;��ұ$wQѕ�����B�)�u��]�6�L���hf�QSg2a�J-���e�G���_B|E�xd��vZ�A�.H��ߓ�.����w�&0,ԇ���ž��4�vΝ²vgl�$+�gI��Cd�x���������o�e�m9�$��a(��u��g��	Y8��&T��%�Y]2�1U)UG�nnT�Bg6�ڊB����χ5A<�)��c��J2'>/@��ĎXo&�fX�M�Cj8���������W��)��t)�ۂ��R��irF�=)<bG�£�@c�iK�놙�6M`d�+gaң4fV��o�%E'���R�*��m��?G�q8,[�6��p������Ż�Ŭ�;L
�`8��}��2�#��٘�0⹽�f��յ2�s|*g{�#>��ެ�*�W��h�Mg�=���'�����>`-��xF�7��,�ïd��tf�!�w�N_��i�5R�B�y?Ց�jՐ�r|�Me�2��]j�k����)�'��^��O`l��R�@��%��4���u�~�D����x�u�"׊@���\h��t�&���w�D~/�pW(ت�@����>��:�u���߮M��fT��Q|Ǘ�)\;�5�\2�b��-�,O�W�3��B�j�Э���8p� F��H]���t� o�!r���s��,j�3�e�)\�Z�\�"v��Ӯ;P}*�%�r�P�Hwc9��gȦd�*�D^��H�l[5�@J7:�a8\�5�Ǟ�9����0o:3��\O�Sfcn���n4~�x&�^���/�[��8�S�ܜ�:ɢ&a킊i�%ϼB3L_+��y�
���15o݈�o;�����պ�H�x7����d���	��ٸcq��&�O4h4G	C(�$ �S�P�I�\{W��?�.SX��
�� ���EqPpd���Z}����LnX��*�1[p6A浔�1
�>z_�o�*�� f�dUꏔP4�;E�=�[a��-/3#�����sg�ū/K�������7�����WkS/��h�#ۏ�^��w*~t��K����a����%�(l���[��G!K������9�'n�l�7�"��}�d��c�U�>͇�s��%��a&"�k�J�wZ��tt�E�S�����2���i��"�k����D��	��q�rE�����H��;00��F��Na�����R-A�7e��Ӹ#h��;):Ԩ��b�\�3Ϳ�)r;
�.�0�~Xiڷ*���I:[