XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���PJ]l��V��b`M�.?�<�e�0�;�<���Õ��+N1Cs�{Y-����ߎH�E��|v`Ｕ�]0`6����Z1��j���Mu��d�"ȷ�t�lT�w13X��|�s�3gb�0zֿ����yp��m$�Ai����+\j�R�rF�4�4)�J�.r�1(lf�,)�`��~����es���	��(��l����1)�ߏ�(��ڦ�k]�/��H�F�O�q�RE��JQ�Z�Y� ��+�r�X�}:$fl�49���_�n�T�t�Bפï{��ƒI�)�=�/S�͚�:�%|E��V�q�D�Bo����	G�����}?�z��w�|#=y������v�u;~9���!�Ơx�	�]M�0G���Ğٌy�����
�aiIƎPn�k�ˀ�*g(s?��~���3|g���t����N)Q���~졕Jr�I��u���P���}�`ram���E �fi����(,��,�n)¬E��Of�=��>ݿ71)|Iu�>f��QU�/=�:�_]��ٸ��[*�y� 9k��K@��!��^}XhP�z��D��ה�E?�]cƨz���5���(G+B[tQ]�_��%�˃ �+_d���/�n�7�@7v&�R�0$�N^ϵ�$�XiG
��(�1��j\�"��YԚ������
sId\���&��b�\��nT�Ef;E���G&���CK. �B���V�+�#V�7�dC��@B�8Ko(YŐ�]Ϙ����[���4��CXlxVHYEB    6867    11501�9@{�9�W|�$~6e���tF]g����"G�).�q�Pu��F��a$R%�qh|-�5	T�&:O�ƺe]Kpyώ����\�ǹ#��0�LPX��������o�}�Bh �\UB��"�VA����j�Ρ��ٿ�<4���jyf���E+q��p\H�PJ`��t���pJ��k����<��*��c^>=~ݣ�~3:N��B@�����)}B�
)�n��z;�>�x-��jG���_�f������@[xC�22�[<�A ԘϲYU$�L��+�M?���
���w��u�C��
tD�=�}�Iy,�W����t�X��,�heI*��
���Nq(�q�*�t��eՍ:���iv���vgj�@��>�Ntj�p�8������x4E�nJ{ �k���͍�����8�K��n#ƫ��KmVk��?���r�~�4.�Rr�ူOᜋ�"?d�;�>K�����_q�(���sN�������f^F*�fM����n�ά�w���AR巭T8i���QIN�o�� �#�U�ý��ʾf"L8����	��m��ao��p�~)VA4'q�+D&i;J<��X���+� �"��zHD�{�7�S!�5�C�}h�j��)�~r�i�vs�s��ץQk��(��Z9���jB,o7᳁����j�y�-~
fUv�م8�mP�{qAV�'�b���]�A1֓�9����{�%.�����	�h�DË�m�b|Iez��ҫS�Z�tPJ0W$��U��+uxFn7@h	�~�tp�������!ӵ��Ի���斶�$ojr�p{��3e�sA�6�"�>%	
������k�$C]mX	��ۉ�����U�їY)�q�����&,�&�V��F��� ���ެ��L=RO�v���:�M�"���}�����p�)��_`X|h������b�#Z;���UC���8{����DXr&rS���7[��q2��=�$KP��+�/8U��g%ci?��?�!����r_pV`S�髆Tj59u)m[�GHY�0��"Rb&M@풷H�ԥ��ļ�}I����eJB�ϐZ@��CI�ۧ�3�&g4��֣�<(�?{��P�$�� �j���E�7�U�%��b�^���,&��-�f�w)T���b�]�SR�Q��ciN�X?.���uUk��,��P=Tt�Jҵ��!�N��M��Wfe�9���aMQ܈���9�GF�FV0W�b\�)Fw$��<�G�kZI�RD3����@�B��<O	��!B�V��e�n ��?$ngD���$N�69���F1B��b�`t1p.�J/f�M�q��|8z �*[�����F��~٥�N<% G[��j���7��-�=�ҏ;��&���E��/0 &��$�;�[ג�1֟ݾ�ggT�(]����{��m��O�kM����A�!]��J/E*��!�]��~�8�2�~������3vT5m?p�7x�X�o�&)3�ALn'K$�Kȝ�q��2O~�;V^F��D�S�q@ 6H�ygڒ��	\&����:�÷�U�^�X�y޾[s�*�𐋗����4\��)�e��������+n-��h�q)�'q�K��~E齛5PW���,i�\�`�])��F?ܬ����Pg���ׄ�b��J���`�� R��'/~������Y2Y��o�/CTV�Ҿ;�gK6�@�[~�i�9)��뿗����\Ha��u!�DKr���h�͹F+""�O`n�{H�5p�	�1F.h:u���ɇ�G�?Ȏ� ���,�]2Sw��yDx(Kj�*�$y�@�i�q��d�5�&�� �`�C@����b_���$E�!UD�!����f��٫L^3,͝�vm��L��Y��i|kϦܐgI���P���	���ҹ4,|�]z5��8��=�N|*�\��M�赕��:1!����3�M7$C�f�Ɨ������s�"<5����'�3��V�a�OǞ��w)}x��fx.�Ї?�S�g���Rұ�mH��Q��r5nS��I��� ��;�%��NDw��d��]�� �i��yΚ���+����������o>�d�F2�l�2S;&
���3^t����ul�K &����,'ԉDʹS�&���������XQ���i�Z�d�s.	H�fw��Z%���%S�TJT\���v��qk^fYS8R!�D�j��=��`X��c��#��6�ˁq��NG�ɑ\V��'h������G�56Z�7`-������?WK:�[c���jǒ�]�~��}�ߜ�I���8+�1�{[����.����?$;��{�+��Y6�����Fj������wfڅ����֚>��|۲m��d��Ǟ��2�ET� pF���ц[1�KY֟���1�Y' �K?�,f��LfV�S��DȢ�%�2��"��3a��s$ws�qs1�ߒ�:�:対g�IȜ})��,P���T�@���gZR���W�q5�[��Y{�?Ȱ@�_1?��B���.)	d�)9ځ����yO2/׹� �t���F��<-���������T�=t�@G�Y����L�I����.<��}�	BW�n2{��L�Q �����B*Px�qm��@�,#�Ҿ���r�s%���dw����!�`��n�J��I� C�XX���$]�'�J��ՈDYG����}�Z��'��cZ�*���iUcͼ>5��ݕ�[��-�X�~�X�A3�����K�m7ݻN[��Y�W��g� �O�׌�y>�<��M�1���i���K%�/o3��Ek��9n��t@t�ÿ�|�;J��}g��s'�I�����93HM��6U0���괵�ױ����\�y�J��~�L��=q߮��õcꅟ�kc"WEW&���	����d��f� ����|�F�7:1wr����ԧ�J���v�WR�bh �+l� 2C�8�p��'Nz@�Wl���+�F���Qp�[7p������2�w��b(~P\$g�92�sBcW i�c�yI��,vC{Q^py_�g�BRc`tn3#@���� �h�jO��o�='4�o�ʇti�!k��k��I]�����޲�ŖU�F�oh�/�����뱧>�f�+�A�V,zx27�5�4 K�U ����3���q9��gv�q�.a
�>B���L/�����ccY��f�}�4���H%.v z8x��@�oȃ)����C/\��� Ye��7�l�Ͳh�^?0;:ZO������n%��DZ��;��d�0w��~X��棭��'y���GD�9�֘��k�xQy�޺��T�?~ �1�zJߚ���yU�ԊgT?�n�ɉM��f� q��qX6^z����e�1�sM��_D/������#�������G$��#��N	=��7��egp�y n�LK|퉹����qb�o""ҙ��]D�0�s����1(�a��8 �Y$�H��~z�4��R��p6k9��,
�E�D�^>i �y�02�fN��;��u�Y�5H��ж�0<�T2���x�a�˧L��)D��,�!�9Fzs7^�b�� !:S�s��!�,E˪gF�=���o+��-'7���o�e/�<�<�B��"C�(<���*��g��3�]H�
��H�)��c�����A�h)���� ��EY�^V��NK"��Whi,'�K��L*��)���� -�[�b`�aqdop���ń$�c�շ^�nӗ��������~�� ,�s��M)�ޑ�~"��+ͪl��vE�ui��h��e���τ�
4�u�ɋ��ϧ��Ħso$p���μV����/�A��s��@��ܢ��ILO�^3/��~F`#C��b�x���]����s��� �ظ�\����EY��t�7��\�Tߍ�@�d�K�J2~�A����:R@S_{�'3W��ln��_�~�%aϘ�b���0�<9���`�|�M|��z߅+��N�[�X��@%������"m�@����,�ԑ���]�E�j+H�`�1��0��PY��$��+�%�)*�	Lb�}���T�r;�;�M���} `�cmȾ�e"y�h�=zz��9�x~)� ����\!o��vN��@SG���y�h��z]���IFr�C*�&��I�)!�͠$"z�;���B�ǀ������z�����52"���бS��s�g�X�5R�Q�'��@]�TSW%���%/��>[�n Y�dG�B��*�p��9��+�h�}������.4���Ղ��k��\j�57��t�3g�eڷL��A�uJV�����$g䞗�	�=2 ?��f��D�Byf�l���b���NF�L�����![l���M��ҟB�WIV'�oA��W�园�B�