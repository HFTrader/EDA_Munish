XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���rc���/}���)6rQ���!9�^��_ʗ�]V~ej���oWŪ޿7��y�r�ʏ�xo��ť�WY����@�`�������g&�5q���nf�k|@���D�5����I&q"���w��4�3u��g���8ұ�j0��i*jR��P�:P0�5�N��G�\�����(��+�/�3���Ĩۡ�!<<)�n7��[�̧��f���}֓Q� �єO����Qah��܋�X\j���������n�F�猫����nP�Nث�	�'[�π�p�K���*&�Y+�#�Ӻ��%$����T�5��kB���xd�&��DƔr/<"��������ZE��� �EקF���?�3���fF����DY�<��+e��V�GnI���m`��bd��,� �2�o�B��j��q6�.�!��$<�ݽ����~��+�? ̅u4�zZ\~N�q�M�_5/�S�T��|��\UAH) ���J��t#l,�D>~T���vy�a)DжUH�M�A���U3pp?�0���^*w��R͓�/�ԃ�fWA�\/L�*��Ja\�<�6��r]��Y��3,¸����)+�a�xh�R%B���ڔ�S#[dj5�h������4(\��{-u�偈��5iL����P�p�&���Jf7�L$���S��߶u���?�TC�^��{���`�2n��*��CP�QIĔ�o
*y�x����z��Zti�c���dXlxVHYEB     f7d     6b0���2|Ɵ�\(Q���쌥��҄��r�o�)[b^?-�ӻ��;���~�
E��!W\1�O��2:������C�����{��G��ʻ�Z���yh��66%�I�b���	! �2�$ly
�YR���i���N �,�6�vW8KU*�N�zv��wZ&��6?Q�����ѳ�Y�pʊ7|C�<��L���S����?�x1`Nf"GƑ^��~�{�&E��?�j���Δ%o��?�P�
)
����� ���!5s]U�A��|*h#����@�9�����$�|MY���jk�kb�_�YJ^y�ZC;�I�߳���v��R��"��lz,%6�E���L�������
4j�=��	�W!�~�Ķވ`ك����qiY
� A]C�_��"ދ;�`^�j(�M�)��9��%��ݞ|)]9��O����!���b@x����N���n�"1܉�����i��=�	�``�f�
\T�	�-\c�{\ҐQ��8~N���TE�A@#6��W�W ��mu��&����¿�2֤r�o?�l6��[���ڎ�(�~<�\���ԑ�uٍ����8)7x�BO�2��bw,����@9Nےs�~�����.�:���:Up\��Vf=�C����?<ٷ|H��@��V���q�4���<���#5�-������&�"�i������)WCRRěeş3w\�ۅ�n�R(ԢOSӿJ=�=m�x�4W,�m.����C��R���̑���u諡B���ѣ�����yD�h�/��8"8`�8@�ޛ��lslϛ��?o����I��8�4�J�������{�*�q�d�pt�����9��q	w���HB�M���������4p>0q��k�fh����6�ݓv��T��H�&��d�¾2E�<%���,�h���G���fj���-�Nf��z-��<�|��C+ڊ=� ����!�]1\a� O�^�[9T����>��I��ʧrׂI�R�1tv9~�z?8�	!�?�:�B��g���/$�qu4`�`�eĜ6�)u�!�Y�R]H2eѹd�?�e$6`�:#-W	�K0D\wv%�nVR��|%b��{��%'��-Ij��r�H��ߺ/��8�S\���N0��o$�.ԁ������K�"3P΋3Y�S��k��T��W�"�܈� ,��z�L��,��;4WY�U��Q��/q>:�v'Y	W�etV\���5�����">��x-6�i���"q��P�R����ZRj���Y�%�\ѕJ� ����e���SS�3�L���c�r`y����0��|��?�=�N�x�i���ƙ�@�BB�>|2�� ���.5fP� y�T�|8��+�h%;����_��	�^Wt4��p��ZIG�Z�)�F'g�:�6	��WG:��/�'��e��ј� Ȅ�4��_��Cql��;�4?B@�mz�|p�7��wGt>�j�p��N���APa�u傛"rrZg\�/��޲�@k�I�4sJ����,�SA����>��g!���s��[v��eZ+T�X�S��+5�t�+�w��P�ࢂ4rDz=ڍ����s���l[��R5}_�+�[\��*Y�;ЦF_l�"��^-�a�6t,�*rH����]�c�:���R�IFuȸ��y�^����{M��