XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=ϴ�Қw>Du���H��!8����4C2��d�]_�C�	LN_b��k��	*a�ZY�' M�3��w�����Ў���G�]�S.|}��@�?�0�J߂�$�`i�cD=�	�a]wɉ�4�A�5��g�0�P�+IOF��2�"a�6���0Hû �o�~k%T�Wœn�,�^�
=��� �D�R�����c��,��ޫrM��<�J����?Q�p����K%����E��|�q8��f~�&4]|y��УW�S���aY7�w�]�%��e��eX�e����5�7E|��8<@�a��g�"�����ⶣ��z���5U�Ȏ�X�D^JU��7�J��Bnlc��\�pK��c;�t_	6{�:^s���¹�ˀu h�-.'E{Ŋ�}�i�I5=��RY� ��y�ƭl���޾��T|�b��Rz�F���rȹ�n5|4yvm`L�y3�q�7�@)����ߡd@G��P�v&�Wq�B��P����j��- $z8�îb v��7�Z$��5���ٙ��8�ci�}��ȝ  ����6�Hf�e��nNRS������/]���O������UyG�3��2�е-1����M��t*j.]�	C�����a�xM!�
d�6�K���Yt�m�p<y��k�b:[`9���R�����������·���F�JSwZ��XBӮ�^"2N��A�(ˋ\��B� �PNG1�-��q��}�1�*ũqChV��B0&M�A\np�N��<��{�:(���Y��ҶfXlxVHYEB    3927     fc0�B#C˫%��@�eX�ǳ�Z3�����g�G��g��0j����k���ϸ����eTD�7������Z�7/eߔU��"�h�:k�_�,+;0qˤ�"B�I2�9��3'����"6:7�!2�A`	+!_2 �/2�p�NsQC�+�6�Yd*y@ͫ��E[T��kT
�Bsz~�N�M�|��f��l2����0�}����d��WK�t��������k]	y��
�S����haЇP�o�g���Ճ�r2��u�����Q�$5����Ѧ6��:��n��ٹ�:_��h�pŏEG]��8��,1�����"r��ړ�d�9
�IK�L���I�P?�����t��\6 #�Oc���7m۩Л
��IM*�	.��*>����|�Y:$�_&'�í�B:���`oݖ�=�u���%���⮽��S�N/��j?��IQt���zK$���q�E�d�(y����k
B���򠾣a����I7;8�'|�n�tG�F�<��	���|���9�����jqQ磯p��~�E�Ly�+L
�y�fbw�9�q�s��j!�k�Ⱥ���@>eTHʠQNK���K$��(h*�E��?�z�:!x�uy�!\?B0���zg��W��R@I���Ã8��fGХ��̴J����mU��>!Ā�Q���69h:H}�Y�!8S7j���D���rUZ8�\3N"poK���&����_�֙�� ���<Ӳz��"µ��K��d>�h��n�b�pq��~�����u���!H�}�o�w�C��YG�\��(Z�_c�Qp]ű*~��T��g/���	+����Ğlb���b
�� D�zS9A���Tr�����'����chO���z��C��1��v�CS��U��Ë�C���ۣ{;�݋M0�	 M}������u�I�g�uK�q+���	���t9�6a��B�vi#��|0�mԥ�٣M'v�;aB�m ͙C��]�闩���H����������1�u��j/�+j��fsn!�� \� �H�b}�p���Q��]e�>i�t�tC��T�I�FO3@��j2���Ӏu3H�M&���b^{����Q���#�In��/�?�N�6x��|&�-~z��O�NgX@�x�ߊgd�)�%�o�J��;����U�H`Z��̅��w�p�>���F�7/�Aa��A�.ߡ����U���먆T&�=b�!Sp�V�6ս�{��.�a<{�ɽ�H��d<V�;�l�RCun)y-(�s�(0��X���<��7������Cp=\^����-.��6�\bP2%k���4�Z���� ���O��!Yxא@؄�DL��b���v���BM�^S��q�8/_r�Ko5pbs	�GO���B������} vM���?��n� �;�.[+K���&�I
PvN��/�E?�#�ԝ�ԫ��	����|ݓ�Y?�u@�ӟ��G�W!���
�T�-��1�=(�8�ܧ�S���D*���P���i�8���p��g���ى$V�9�����&��؍@�)��>�̦�ً��S��cUD�/��>�u�������^��G����`3��������ˈitk'���)1�|Ft6,�ؘys�!9��m��q�k�¡q�1���b���sw���mμ+�Ľv�E$M�ٯ����)�5v�m��.�R���)��QϘ��zi����tҩ��A	H���oX\|l}��w�'s1p�9F�,2�C���e�ПH�I��ă��¶S�<�1/.��҂v���4�1��鬫�L�@ҭ���	/����{��}��#5Cb�;���­�/�l�\yg�|��=Wb��ݻ�qO Ci�%�'�y�k��N? ��;�|)4���,�|O3���IH�!�;d�w�Urs�XF��� �(uL`9U_ëR�d/ˠ���gf�U��r׫�2>��@l�)r�8Y�tĭ���^ b\�o~ђ{k�_K&�Eކ���ȳ��S�&#��a��1��r4N����OO�^6l�A�~}�܈���7��j��s�8?�E:@�i6��v�������SԮ#���� �c#��Gwyqt�>�!1������sݎ�]�.6�u�E�
?�֍@��Ϳ���Q�����޲B���@�4��&�E��O>?� ��R(���H=�h�O�Y�@V�Yu�����j���/��7��r��ӡJ$�K:���7���2! �/�`T=��ؾ_�	�>�X	��R-Ɗ����
?[���. �W������-�0Dj�2&��􅫛Ǒ!Yu�2L�|��^�	u�RV���-c������������z�.��!�sA*=�Q$�S������4m>S�M�� Uϡs_���
׼�Wzy]��y�gD�XʎO�\�#>Y(]��	v�X��h��`ʰ�$�IY����쉖��L["]��&��aoDcdY���.��!���S�.���Ϭ}QG
�Ȯz[�c � �cY����sGh1���H�K#KF�eC�܅�f�t�m L�f��AZ�8Hn�R�|�:�� j�6mi\���93B*Us�G��:�6;��ϴҽ��B��L3+�J	�$v��
U�;�b��#Uu�����|����J
T�6so��*7).X��,���Y�#`��L����_������c��E�7b�KH������}�x�z��o�)�ZG������?�5�`}�s�;t�I>�o0ݖ��Hd`X
G:�OP��g��F�$� -^�{j x���R ���r�X�j��Z9VTZ��z��w8��A�E�,�н��_t�$9�|ow�=o(�JW�n]&w�~�n��;#��kCY�ȃ��B}.�ڔ�w3�Wws��`�Q�]佁���O*H�v�Rt�Y$F�!X6S����(�?\	����̩Jl�ɤ[��;��vH)2����Rb�<��nȚ$�����{,|���G��4H<�pN���-�ι�8h<����+��p$������n����b�i��W��K�5b�w$x?Xw��#��1Y�qV�S�w���������[Ą�)�}���TZF�����V�Z�O�Y�u7Rn��%�5x.�'���R��Ե�~y�01�%��S�Y\s�w;M3��~`�����T��!>��cޗ�XoB�pN����L� )mr�'��\�����ϣ��;G�PbL�ZM�-�s������}QR5cn�H۷"�z��	j�^X}����k�<q�=�#[�2��!�Yg���� �>��2G(OP��>�7+�J���-.2���|=QE�K7�"��Dp�%��.�M�pܐ�����ρ�C�c:�d����L���E�oW�!:�p�yw�+s�{��r8Xz��g��Xӭ��O�C�dۙj}��5 ����J��}���[�B��J5d���5�|s���T[S��:f�~rڮL܀ ʷ�#SQ��ҩrOl���R7f����D�<����]��R]�������I~]�@vu7n@�g��%���qlb	�|�dݑ�ͼ�_3e�~Ӎ%O	is\���NI_)qP����
��*:ֶ<C$/����Xyu��U ^�Z{r�tr���q���1"�pu�����~>�O��޻�	�����[!y��1���I=.5�ם6~��7Ov^��z��d�m�P��溱�z���b�Z�Ӱᓕ��{�bG��08�Ʈ�A�"WW�'��?��d�oB���3\b�q�1�	�PD;��ן>H")������$"�#L$_�h�K`~�~�!�mE�	~���F��ߟz��N0ñ�n��*luwV�4`(u4�=�0(���K�0�Q���I����g�s�oő�B��'�;S�W�6�Ƹ`�����f84�W �$s��(ʤJ-���m5��ӹ:G�-��Ç"x��C._�G���K����)k��쭋 *ae3�S}�mѨ��<����.	4