XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��iN�@��?ŧ_�!�,��7�Q�A��Z���
V��,|������jȃ�A<�AXG��ש�X*H3���.�v/_ ��h�wq�:Yf<G����pt����%&�iѺ'�7�
1p<�A�M�ySh����c��lK>�����km�b���ܑ"�࿤H�nVdٱ��f�����L,��~\q�,�ɡ��bexsO��G����k}�;պ~�H���°��6��H.����~M/l�^���ߒ%i���:�-�h��,j����H�4�jA�m�j�B���G�3�� %zF4��65�y?k�MQLlY=�-�"��z�m������|禺{z��=~:��~��.�bd�/���o��pgK��LQضE8��"QTI��H��e�V�����	�mw�;6�9h@���� �cS��h��!��M�y"ַR�8�o�R��-�����Ȅ6W$����(�W�C�a~�t0}���*@��2�O�&G03UJ��t�C!K}-o��|��>aë�>�VB�%�1��YO*��pz�d�Q�>����u��z���П�*%H���lz�E����\1
�Ǒ�<f8l���HيR�S`���k��p��6۳?H�5��l#�M�f�v8&�3�� )%�G'�g�B�w�E)_�+���@hߤ���zm߉3��!�D,ict��^M���W�Z��&�����5���SK&�춯�^��3�H�'(XlxVHYEB    1853     8104j�sg��x��#�;d�+��k/���n&AgeQlBFW���v�����hк�@�
5�02_��&�>��i�ޓ�/��hU��SZ,�z��ϜA���c�{��e{�6�pz�L�/D3����Q��I��H7���*�Dg�q���t\�|Lxs���д�v���t��h��}�O>$&㇏�k��R���s<��*��ʸW�Չ���(~�Z!��ݵ�tb������3n�o�Pyf�^xٹ��)N�!J'g�j ��M�¹����.���<NB*v�'�ؤ�&ɲ�ҥjtZOSO�|Z�hL	��^��f��H�r����_�.`���3PI������ b��~S�zw��ey�	�_�Ryjx������A:����H�=Х;��(i�\���3 �2Q��!��T�8tԱ�E-O�EaE�H~�	~�H����o�9��YY�Y���ޫBi�%AQ|�_�I�%Ax�Z��礱t�G�Z4Wa�F�h<����k�^{�	�1�-�wW�]�>6�<В� Z�����ܵ85)�����d�@�t�31�4�Y
�tV���E�XV	���;�:qZ��<^Y���&��"x�~fO$��v�I�/i�-��c����cD��q�|�[I���o� �c��$8�����H� :��T�x�B"��9!T�5 r(���;��p?%s�Gk�%4��_�k�~��hf$|���9x�_���lh�v]j�#c�K�X"6���Od�����74טjyU!�i���{ErOJ1p��먜*�O�c�Jh��tXG̮��#.%��s��%;���5���aCK���^b`Vӭ���]Y�c�xoF���Ͱ&��fpR�JM�Y����ȅ R%��G-�(bzG��#GJ�m�̃L���	,��:���*�9�M�f��2f~�=�	�]���`�n"��m��4M��qrUK��NOIo[Y�d��\��;�C�@�h�Ň�BH5�m�F�Kh��G����M:��	�h��:���p�Z�׮  �i���s����~��ZZz$`|��3��ǀ3HP)d�*g�ʙWS���TJ8P]������2_��y�sW�L�1`V���� 1��(Yȭ��=�'wM��1�-�re�vl��uy`F���c/|�U���5�%�Ν3�,TQ"��.�r�%��b^|��{,�*�4
��^�X���������R���^���8pg7�ވ���zvIbSM	�: 9XG��n�L�[���k�������7����J&\Ů��+��*�;�Ԫ��>zT�\��M>RWB[w��S��HԪP'׋�'Iۓ^��At"6��w@� ��?�:�H-��䒞f��T���~8���h����.��d�����z�yؾ+{kE���;�{sOt�����#�j!8l�.j8�/*b)�5��_4݃�X��8� �DX���J�Lg�-�+�0XM�
$��@<RsI+n�[�����b��ty����I +�M�d��`���U�(��˩c�b�g��sD�25�٨�k��8�h����ث!<Z�ބ��Ł�Il3�Ps;dY���7��`��ecr��ċ��q��ޘ6�A�B
&��
�SZTs����#��(�P�=�����V�4ro��(<\���A��'�,a>���'��fSDs����.��FF��'�!Мo�'7�C �+�5�*ڹi��w$w�(LU���e�A�Ʒ_����/�=PAE�7�[��?oO\��������?.�_�!jwW���n��9����35��%�֔�u���(:ak�M���c��V���G��`?�gS���b�3뿒9&(=~���"ۮA8s�9b &�\Z4q��%&���6��Kϒ(��V��ieVP=t6�:�n(�A'hDu��kM$$4���|�[N4��C��:1w��DϲCW�'r4��L�NMŶU��4�i��	�G���f��#{MoDK$����[���|!w�u�%��%�
�]1�l�,���Eq���؊�6HX�_v���N/�t9gd�ϝ.�K���u