XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����#�5�k��*��2����%/DQ,^Y���TR����T��}׮u9�+?��>��z�S�T}���l	�X7xM_�X��g��"�r���
��V�1�2	p����[*GH�x*_%f�����u�A	�uQ�. 
f\��;�P2���o�T�� 
�GY|H��X���r4�b�Y  �E����"p�����{�T��)���ۨ2�\D��gP����v����qdC����m�2��_�{�~�|7�za�@^u��Upz�>��#`��y����,PMO��5�C�s�{便>9�����m�FY�9Q���~$Ut�`Z��y|<��čw�j���*:���pN��0f��G?�9Zn��Q�i$��V�d=\�)2�~���0��.���5�8�y�m��U΋�����
��Q�����6^m9����m�}-�I�7h@_���8Ӥ�=n�G��&�T:2n`��ajVp7�q��sLBaa��&.m�≹&7�j4�}1�?�B ��HO�ç{L��v����?��[AD.*�`P�k$�� A��$9�Z]W0m��Y�3W	0��OJ���:,_)c%a�����@=�7�U��$��ӽ�R*�6݋K8�%Z���f�i����b,=폪-R5��`?�8�{�`���$c�eb˹'�-�����Ѳ�,��beT���c��#���]�X��S���o�������!�<S�5�[���x�yٿ6;��[�>^�OD˟�z,pXlxVHYEB    1e9e     910�zߕ�9K\ЮJrh %�ea&x-z�oh������#�
�ɬ���y�qoC�Z[�G�&�nv�c4���%qӮs9���&�.l���]�5�����R���Դ��	�;ݔT�hFm��,X
�5A���ߧ��ڞ��ܺ\r ;�{<��C�%ax���;�!E�X�9���"
v�t����֌�����0��j�H~��y۠*-��/l�v��#f'$�m��R����T�x��%�U�����c��"#lic:<s ���T�ד|��wa��`�#�8O�'�Վ YM���5��B 1'9Q�u��[2i��0�h*��IB/�r��R�C	�\}�[Юp&�� Q�5��к�	����M�9��jD��ѓE���� ��R��޹�hޓ�ЂZ��MP�Ƌ�`|�l�H��b��u\�-�p�2v�sC��f
-+#-��C�,��4�n~�?�
�)��c�Ι �4¬6oo.���)�8D�(VjϡSa7�YJ�v��:`LM�}+�r��i��p������T���e������`K���~�
�����W����`j�J�>����m�5O[M<\�w"����e�۴��{mt@��%�$�gx��U��R���
�N���fG���P�g!sМ&�ĻA�@1g��1�Q�����IE����/iщ��n�~�|d4���;c�Q��P�I����N�LTd×��"�z�Ҫ�ݢ���&a��ZA�}�=:�^�X����9���L�Lzd�z�R�������F�̽'3�f�gb�-�Ofq8��`�Q���L8�@�)����gW=�5��� ̈́�+Dl�EGZ�BT�6�\���"�7\,f��{G����&�[�l�OD��.p�p��i
*N�p.ۀ��J
��)����!�-Qɧ�S}������%��B�S�}�2j����:g��,6$y5��`�e;�<�Ŷ���	���Fw�ܗ�=�s4+�ST�#�&�T2���$:z�r~���P����":]U<�S��w�G���l�rw�2�k(?���Š�K�1T��r�#X��١���+Ը��ET�@�A��r|��3r�/�=����2�N�G���Fsj�s�F@7j�ݷ��M*��͢�g�8d�I�q�zD.q�<Ö&j�^�pZ�ʁ�KV�~���=!܋T����M]OA����1݉�74��Ng=ߢ]��N@��;�&u�����q�tݬ&��J� "�_f���c�e?�A���־>��0N�@��tb�srHk��/����҄�Sw�}N2i��.����̗�{��W�p�<%Ԋ������@����|P��O�"�D���#�t-ҟ�+Q�M|��;�*p�n�/�G��{��&/�Me�'�pz���Q[����=����H�d���1]����&W�Eu2M2 �%-�؊�wOb�]D}U)QE˞������F�D��YK��M����AE�te�hx��Y���z��ͦ���==B�~W#��`�K�$F�����R�Ed��,�K���`[9n�_S�Ls�޹27�3}�]��-y�`_��y[�J�Ѧm��p�
��!c�t�4=]U����G�N�o?P-Κ�VxG�����,Fz���+�۹3?oG��/nj��EH�bi�TTh��M��6�=���pIjq�$#�8�_M��}¢]�4˒	ܞυJ�83���Z ׯ*�@ڧ?U�/�?ć�|�[s�X7u�¯���P���k.RO���Y�������XXX��.O��� �`��#^��U���x���b��iܧY�����>����.���� WV��5����Ng�h��FX��ϩ���(�h�y����C��f{R��ro΄~;j�F](�/���y�R�$-����?H㫐���΄���mFfP�i�
��Ij�;W�;��a%I���f�>N�1��)A�K1)d4Eۏ5y#82\�J�ή�mƒ�`r�#1g�a�>X�
P�c�讗��!)	"Z���e����T�ׂ)H�E����w]���Vj� �����h���_<4��L�1{�kc]?u��P�Wѧ1᳡C1��O�sֿ��b�z�cQ����P�����@�T�r��FK�a� ZH@�O�g��	A�w��qr�F$��ٝ�+�E@z�>S��b�3b7����C�kID[쳴U	��b)A�-�j���l|]��������!�|'Bc8\�ܖ{7��r���$#����!�G�U��n%����#�7^�7BG�:|"�n1?�Xz���