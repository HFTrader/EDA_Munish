XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5�hn֐�)�_]���3���9x���	I򦀃�px�w���熄b�-N���=�Z��ݡ�Z���\�H�$Ba���Q���}N�������Dο�ӻ����g���+N�)��(r_|pS��W�(���<�HWR�e;�຦}�������=s���7��c�|�fN�(
��e>e�r�Y��)㟑䠣D/��j�G���r�H  A�v��2^�Q��}��}���4������ĩ���lm�o:�MV�b��-��+A��Q�$*3�Ǣ�ݣ���a��+�n�@j�j�[�J���xW,�)�]q㰘�W���F�0�;,�I�sΙ��u1/pS%.��<�G*.�P
��(�,f ?N@q���Te���&���d�[1WXP��K���$@�R���<;��e��m*�kW'&֯Lf[��̋47��ͅi�~��>m5u
�6�U�n�'slg���,8~H`�nD~�Z�ٌX��'�K��&�5���5��O�Lm�K���:*���D���qՏ�M@6P��6���ф�+�fȃ�PTf��v�H<Y�6�֣�S+6q0T�qQ����66����) �T��Jmm����W�ǣC�Mǫ]�?�D k���lK��2ܠ�^�#�r�5�H�h̝�e���spU�;r��R���9�Ӗ��]�U=����v��~Z����c�S07�#� 3����m�\�W�������u���J��ʴ�*\�� ���rR�P�l1�r�?�q\XlxVHYEB    2f9f     c60m�H�L�*�a� �,�E2p�ը`��g������%�6���<�'���O����b�HVT�5+�_ b��i}m�Ѻ����[:dR�]�*��Ɯ���h�z�����J�*U�eA��[��.��{�x���|���(7p*�as��u(p.</�
�`8��բҷ���1��܇�8#y���7ē�vA��T6�1�9�r�8����U�0��gw��mׂp�?��@���"����a�cnQ�E">h�M#W:û>��.����+;-$�쀶���b8$}�1��U9�N��LXjT��֖�o=�8��g!-���{chx�C� x$�.�]zxOW�֒*��:qY7�Bg�6[���ԡXk��k�J?Q�����>w�M��MC�8CH� � ��h���DPCڌ��AL6�-�3���e���8
�򄒭G6u�*��E@�,�F��@����;,�2�9^>��%�/ᮟ�  *:�C�	��ٙ����"�-��j��}�8+�"4�x�5��@��Bl�b��Z�S��{=e��&�]��zCI���I�k9/71V*;�9.�9�����z�6M�I}���@����(,���܏�ܜ�]6�;���U+��;�U��E2���c�x��khs�%ڏ�hsV�Z����"MA�G���ٻ+�Dv�u�ě�7g�Y�wF�Dl9J�gv�������f��[�m��R�S:(�۽���/�N�x%v�ٲ$D���h����G�����@�`_yA��'�q��~��o�#&:�&�U@�eQK6ng3�MO�5�jK9�Yp�obW����@�e�}@M� �{h;�2�m�!0���<K�0z�2ՠ����  N&ghJ��c��hJ0L0O?1U�$4�, /�7����!?���_��+�7�"�?e����	�������ɘ�i�3��e��i�H*=��p����M�=¿Y�o�?�;�u��г���h+]�Hf��}�2��ju�N���V%�>�'����>3?P%�I\2$Z�zh�� �����C��f��
�NJ��c�~̷ �������TpQ'㟋������ 0�|��
\��bD��=0��,/�B�>"�t��x~&�kD>u#����,lȥ�v�x?��	��UMmi��׸��yd�F��ɪ^�#au^��FF�.x�>��u�ޘ;�hZ��
FR���@R��v��1��ϓ�&�<��+h������N>3�	��P9�7\�Fo� ��*w�+��Sv���K��J�朧k�{�FX���Pxd͈�A���R� �Y+O�K�h�)�w���{&K�#��%��^�/0ZDo�a	�گd��s�s`��tt�ƌzy�kr�c���{�+(�\��xJ�d�҇��ZX���tݏ�F �����^|?58M̟z���D��������s��Z  �|J��v�Wx�y�$��^�!�|?ЧoU5<�΃��&�A��r�X���6?��FPC���T唕��P^�Mw��Ƥo{_jR�,�.iEj��b�p)?M}�M��;�|�'3m@;���z���@~v�T��pe��G�+<�2��U�u�$JϾ}^w+�dJu���fK��FD<����]�}��WS�_1�P7C֞��%�W&��µR���'�?�y��G���<8��B�<���Sy~�톄�c<	ȅ~iAYe����FHݙ~�(}��;I��T���(0m�8��	6�s�.dbv�o�#�rp�x�'�u��_���	!�����,�0t�.�Elt1��^� �����E۹-~K=�@�����Ro�dw����zZ���n��;O#�9�J��%�!����h�C?B��-���.n�ꋛ�=m��Gkf�z���^?o��$��p�F�O)	���83���ZJ��I;��!F�����א]^�R��sA��,��IܴԃQ�zh�l����j_�a`&>)/�GD�H>;X�>��p�shދ'�?<�gd���V�.�D)-�}����ɷ����.x�S��6h��F}�[J�=m�^��Ǝ
_��}�KRڢd;��E5
X��l|��6��_�6h]Vv���:��R����=�
�7��F�*�(����E�u�;�0#�dN�-O9�V�K0	����\
e�WJR�X=ݙ���al�%ĵ���H��k��n�&R�@��`�x�g��a��꩝��/ȜF��b
U��t��0��Ct������`�i�<������`IJ�4?k�"�PIg� �����h݉��H���@�7�hOo���)�8d޹5�G��cr|��i?��d�r��v�G���vZV>V�P�2�!����qr�P�@I䠺>�*�8�G�!:���#�B��ƂZ��^t�ɍR�ҍ�7��K}][D�����0�x��_�fE������k��y'ݒi+�n]`9�}�~�r������F�s=Ⱥ�Z}b�^E�N��Au1�4��%��_cd���T\�p�v���9n=�<����\�"�G�G�$9�'�G�fv�f �|�N�8���*8vF�
xQTVQ�^���)�3Y��C�����x�yøZ#cb�$��{�^�#.�$fכ�`
(��g|�n��K8՝,���W2���u�� n0�ݣ�)TaT-~��X,<�L1;��I�jQ���x(��m����n�\�ٌ�΂��e�j�%�v�����P�Z�K��Mk$7U�[�����Y��<����K�'0���������c�@W\�˚����َ��u� �֒p�&� �@�z�0��;� U�Q+�) ���?��c����I?Q�
���.�%�:WEH:��u������$iE�X�+��U���U{��XL����NU�\��A�?E	u^�����s�N͸��P�I�Q�����\;�� �BkP�'I�O�_%���'��m�Ǚ�fr:>�e!$�/A���վ�Q���nN��32l�iH�P�'
��щ�7)�w����*Q����y��5���D�;/I�;���e����Ņ����3t��l���젚a�yBKY~Q��熷M�ᆳ��y{z�7ϒ^�\8!���5�`D��I�(��p�~MQ