XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����{
Q���EP�8�t�b7�w}�'�W��}�NI[�:U�kx���i;�$&�$d�i�e}ku�:����y������ %�e!ֽ4���)�o}%,_.�:J�\�.�r�yu�%���)�4V%�lz5�e���燄��i7Ň�mD��]���hn�0�8��2</Ԡ8`#x#��z��$�Ek3�y���)��CG>X��N0K�`>W-;��L���T��]Kµ�F4�H�9���c$�k���x�c��l�`v��λč1�?푉�<S��@�>�.���K�Iׄ��'�$7�?M�A�%2�	wjJp��t�&�{4�vx!�s��9Å����i��ONX�"{rV5�D$�B^���j���,�)�P�0K���9��=���sr|q@�ʭ*x��Ʌ�nW{��mQR�r�.�<*�S����G��K��\���!������I��rZ�w�MNn!e]�7,9=?p�����;AÖi����l�HN��(��yڒǋ�s�|�7FYY���.5����.���K�G��6���T��H�><g=e7��\r�u����G�&��QZ�P�k��6�%!Ҡ����s�ë��� ���@��T�6~�	~�E6�;��0�Y
RȌSct+�7x��0�	�n7ا�Η����mg�;��<�p熁D�VH޹�@%�:��4�ëyT�a����(�D��k�D~��/��׎Hm� _ӘB���KJ����k�F�2~�&`߻��XlxVHYEB    5694    1290�ԟ y�F�j�v�0��E�8�k��lG�b��y��B �M��-N�7��&J��
bI���	΍�P
�ъ�s�%�T)$c�G�&�`���2E�"�u��PcS�) Ed���`�{N�E>q�k4p!d�*���6+Q�ً=a6���_���$'�a�xdBrY1Hǻ5�zBׇ�D��I�����D?S��[9� P+��biN�vR'H>���ir�\��!2�ڼ�;�_ZK���tn
�TF���UIM�W�����^d��K>C��}l�r��r���ό
�#�����\N=i�p�:[��V�&6�0�'yVZ*2�lyF�@��d��Y������u�����D1޺�!�O8qҞ�漸�Q�l�����?�ƶ����n5?za��H	;����"C����c�|@�qR�O;��8���������
J$ ����G
�yp2�KM�|�ƽXP�kQd�x馦�	�[���a�*�('QDX�	��*	:��.��Ed�4V�{�SܙT�d=*��<�,7��vJ��u�cB�����+Ni�q�P�t��$�Sn ��F͔<��D���n|U��DZ_� o�"Ӌ��i1��B��<`�/����6p�M��Ь���o�����R��^���^e���h9e�I*�v<[S���¼OÖ�'?G�h|Y;�f�6Xİa�[ׅ��ʶ�'q�?�FM���u� a�G�f��c�Mf����)�X[��ޅ� Z����Z��m��n#��:Rin�e�����ܢ��E*�� 2�VZlu�h�
	3���\w��4V!4�m*�mє��I۝�#� ��o�&0�{@҃]6ek��u
g3�Z�p��N��mv���CԤD@�۱�[���D�I��uA�0��u�w���c��X����#F}�gF�����ζ��,р��֡���x�[�������@B�4�	Is�nI������^U�FCdK椰��&��qe�����b����߫9xA�e:G3_�2��c�L�=�%�H��Ց~ĝ� �>z
����VeS���6�z�H�R���*�1f���eX�*�sk!�=IY	4'鬐��-O�������|h�8�楚^�.Vn5y+��}�t�#{)���ɵzF�nR�F�^�&.�X4D��u���������&o!�蛇�@�d+�b�����&��� ���aFPWf���%�-�x�X<ζm����E�g�]ۇjm�-.��9D�}��> Tvlp��N�Ȇ���Ds��1�G3^��F�s���s֎ Q�wX�B�p�?��������\�qs.��ܖ�%�(�m�V�
6ڱ��K���I~.���iOa�s.~?����N}"cn2MC<Bر��QI}�?��EP&�&�󁃽�=�ljb}�8�G��8�~�A2V��&��|�d��@��RD_�ң>VO�`�N�;4v�?�;�u;AIi@�#2�O�Z'C%6�8��ZP�&-���ƃ�����h�wR�Tq�w�C�ady�	�Np�_l
j.{��;qTP"�6�1n0�R.�DL�&w�{������(_�V�Hr�Zvp/�^p�	'l�<�G��I%�zѷ�U?e��*d��4�4:�^N����p����>r�vc`�q�fm�m�Y�w!=�\�+�L���:Ǝ2 c���A�����8�s�7$�r����b��.��2J(��_����B���Ēϒg�q��CZ�Kh=E2�\��5�yn�Ҳ��d�|��m�`��ߏ��r�v�s���^��ag�z(k������h�� w�k�:(��u�B(�m�@�U�L�6��t��I��L X��'t�I���C�������&�~ah�\=��/�L=��h~��@�Ug�oa�Ah�D��6!�姦KG�1�#r��$0��98�S�w	T���l�y�H����"��Z�.��x>i�-���
�L� G�ki[���2�XZ-�E����L�/���Jz�R�p���p�2�u�ZG���Rʽ��f��2�v]�O�=�k��RSwk�tPS�r��%�b�/�"�/��=�)C���.ݜ���d��X���0�z������Ba%x����C��ߺ䐉&T;�´� �� g�8�l�ғ�,8t��!�ޔß��fNQ�P���h��7#�4��Y�(Ѳ����j܉wԟ�_�͜0y/3/ 
2?����#��i�+f2��o�Gc �{�'Ł�c�ۿ=5Vi�'���?y s�<3�.�j�Y���x���Hl������K��}���Q�IK����A���)�v�{`I�[`�m���Qg��UY8U�}(�����u��$^�Y;Za�+�W��͒��MjQO�iU"T`�>Dח�4{��ǋ2��p��u��Tr�(݋Le�2�_!2G��5��{�K0�f�Y\+MBMI~�`�e��+`�p��p^"Y�'@?0�`�6L����%W\]���U��d���nL���*)�f�~�YG\�_�ZD�m0[{s9@'JY9����đ	����ԟ�H^�"o��ޔ�v�s+�`��ܱZ��A��	�	+�����_���%9+�<�o�R�\�8`���זt�n��y�xU�j���ҋ��$�\�l��ŕ�آ��l;��m�	腟)�EGKe]~Ӓ�9����=�.��\�4���G�s<a��0�Fm�ì?j�j(]!�U_�F�l]�rB���jծ3J?�z�߷1벅1�x�Jպ1�k���u�,����t\�8�ه��I��U��s�D���:�\�Q�!J�Uy!N�EP[t��c)��q��(2�M��f�� u
���R4�K�1wzl!�܁P҈Mh~mJ���Y!�_�����a���gg�${l��I�h�"�֎��]vA��.T�iS���������$&��7��M,�](h��W�FA�gV3�S��MN��򒟟�D���e�X�S�����	R�������֑��C���1��m�{���5�»�z�ΐ ���9���5���#��p�ߒ��K UK�=�e �~M2fLՁ5��N/0m��d����2U�D��JG��	���>�S�Y+Ɍ(���S��t�L����a�_B�{ի�������'0��Dp�f��Jҽn�Y�J��p���ءCч�eDg���usU'���f��V���1��c�p�TiH�Are���Ɍ��Q�<*<��v�����m�ќ�'��LY[rT��&�j5Y�(��i�7l�e��q�BZBP��.�} ���F����T�ţ~���sT���&F�OV^�Od�')v���śJL2��(�������i�>�\ ّ�����b�>Q� O�������N�b�}�|����� ق&�Y> �y=#��"7���o�YXJc�׉6lA�]oG��ـ�np��N��f�0��m�X�Xt�#�$�u���I��6X5n��'�>�R��E�������p����#�b0q�B�4	�9���2���ז��[��Hf�a9R£I�#5���E��n߷䷍"���@7v%yH� ��`��K��Ҁc�O��O��G�Hft�8豣�����Ix�}��c#�MFY�X�/����J(^�T��\r���-��H];<�ȴ������∆�3Alv�S6���e\i�"a���P�-�����A�>���������7ܾ�����|D�2��Y 8�8.iQX05_E�y���H�5�0&b!�	��(Ҿ|
O-��Pͫ�?݀v�P�$��w���g���obʁ	��P�K$*��V[��.�lؕ>Y����^����Pol��l%s��+�8��ٜ�{����i�G�H���?�y��]�͢է(Q5h�����y����(�����W]��m��T��M����A��{JbE��h.|�v��v�o�0NJ�5�o�UtX}}���ո+tw~Q&�H����� v�ak�/�b�E]'Z��O���Ѕ	��%�	Yzxҡ���a'�� ,�L��}�l�^��U�\�qʗj&�E}�[�Y���V ��L��.+/盇�WU<�}��$@�l� �d߸e�b2Z�C]h&)��yhn����n�E�J�<u�¨�� Uۏ�?�/( �K;��q>�CN�8l ?H�8��"���u���$�Ƨ�l��,ם%�3�?�٣Z@�n$�}�DȢ�@��i��WU;�==t�!q��p���	�����@�I<��2Y�ʓ��;����1��"��
zWfq��i���{�.A��N��8�L}�����gTT�l�^��]%�Kr	Et�D�R7KzH�5���� ����e��B�L����E�K[ϢÑ�-5�3*`e/Րu%���c6����J�C��x�~��s�	���4����alu��S�j^�-MSU�s��I2_�p!�~�(@D�:V�i�vJ�p@�`2�4B@7B�R���{���]OD�TH���w��if��VJ�M�S<ŵ�])��K� ��]
"k䳬$�Eb�:
�����耏b�F��,O�̛�a�Z��jmN����Dd�s���hޚ:�L�8�J��v�ʃ�j��m�`�m��)ϛ3"8��*jƛ�s��J�v+?#��Ul��@���eo\Sl�43m=��*̙gƐh	��ޟ)�es�P'��-��5o�4^�:җzƊ9.���5�:|�)����i17�w�0�DD�k