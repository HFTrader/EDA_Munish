XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����i���2��̱��d��S��k���yh
 �Ml��(��6_�	���ӑ;-_~�'T�ļ�V5Z�;����`���,�i��b��va��)#�.��W$A�pF?�o.��LQ^�*�RP	_Z�|3F$�w��lN�]X��r똨ǹp�`q�ǜ�p� �߼K����`3���J12e�c�R2։ K�Fnd�[g(h���.��a�`�՝��N�Z����d�Q�������܆��͌ �m�5��L�<$���57r���)c���˖�������,T����O����G����`_�Ѯ��5�M��-ĺG�7��j�Pt���~&k��-���ХJ"n�퓒��]v'Jt����cO�j���o��݀�_,4��1 �_�)g771�����(�[��t�[�
�q:�>��=�b��U��&�Y�~,p��|��r�r�.qowH��Ƽe�ݚ��R�|�) �i�`Ӱ;���蕏zf�ػ����`˓�ӡ!gÐ��{wj��4,F[ʟ[����ll'��J�0�O��~�G!?�9#�a��d�X���8fB�N�L���->�r�"h_Q0�[�Jd�?��f�8ÅҢӳAC q�p�G�L3Ҷ����R=
1}�B_
W�Ap`�R� !y�����$5X-Y�sq�����Q:g���︎ľ@�I3S5 �x\���~H(�.�Qf9���&���4��Е��ce��k�l>f9#��q�{�Y@`� lhXlxVHYEB    1a5b     890�h<���[���X��&��l�h� v�F)�¬�(]��o8�>�i� "�6&�@1/e+�m��B��B@;�o����M��W��?���f��e�U�Nw�����Q�V�C���er�� "�&�7��g:'w��!	M4�Ї
�������r�0��#�6Kzp�0�ݪ�3Ǳ��5�9�9�Љ��K��ǚ�T\�|��ϊ��c)~��#Ci`}�<�n�ipF�l*{i�FVp7v�sk��$3���-��R��� 
(�'�d�^zJCX�00u��Qs�ܾ^j<Hk��Ix^�펕=���w�-��9�����Ӻ��yT?����편rhW�f�䶘�W����ӭ1��d���M7�z27�3�z3f;1�o,3��#yhk�'��vZ� �D����].�7�W^4�^~�Y��=�&�e�5��@��KC���rwd+z/�Z���jQ�(�ٟ�[�ߝ403������I@˭��2��Nx�yy��O��"�֢ՙ�$D=�G^yVߠ�&}z7�y]��jIb��:��C[�;l�x � N�`�E����sJ67;���8s��*��hq�`;���	��.η���D�H�[Ֆ�[lK�ǆr��ߙ
2F�u���{��4�=��8^�7�I�eLŅ�ˤ��!I��c�ѭ|����M��C�sJX<��KcL���J�]u��b*�S(� ��z`$h��]$�rK娃�YMqm�2��"�!FD�f��%��?"���d��ƭ����8���8��æ7��s��c4i
��ؿ�N¥ڇ~�A yU��Fsx���b�xTݸ��/��``5\�=�����@�[��m�� t�����0����nL�WZ�`��n�B�ꬂ�Y��dư|��@]�����F�"�~6*�5rt�Z$��_4�B���������?	��.В��2;���t%�^��Ua�e��`2�Bi��y&+\'#8{����=�4��A�%Xe�޶�� .�s���'Yu��
�R�V�!i��U�����s�ufqx�/l��Mԑ�!�ƪ O�l�t��׿�aZ�}�j\��BA�J_�<�W�6].s�a"a�Wi�]�tg4� �u�Bm�.k dr�<��[Z��^�/Lb}�� �Pqv1�U{D�ǰT�0���o��%v*3r�Y]=���5�K���U;?]���,�N��g�O����3P��]85�#���ʧ�*-wu#��wj�\�/��B� ؚ>�� �����v5�<BɂO����GDB}$ރ���_��b$u�s��։vxq=���i?�� ���v�3NV����$��	C4�F-�0:��ahk�\n�^��3rC=�yP����y֮m�ϽSq�z]�˘R)c�t���,v/��	�Ϲg�.Ώv��Ǧ��ht[K����f���������4�%�����M���´�!;Xit-��k^2��9X�[���w��S�Vt�-��]�:Q�����C�������w~W��0�G���)�F��[�M�����ǵ���>�[К�	����F��N���F� �ChrTx�`��ݒf��A�@0�8�H�\ZX�2{apC��f��z���ay�b�4�iR���JVCFj�d&Χ]��_!6��I֙�.{�m/�5�x��p:2�8�8��2��Tĳ�����NNQ�g�$B˾���g�)	��&� gf0z���0CSTm��m���z�a�o�A��{�� Zз�#���o!b��)�:�"V�p����S!G��-�H�$&�[�^�,oB�֥�j�g�ٽ��le?p���Ϳ��9���;Ó:�.�*�_gS�,+k�#M6.�($����+qqU�9�3��r�m��q�|�Y^`D<��G���?@���ik�h�������	N�V�����z)�M��M@�T�i0,��\׀uDx�M�Cv��m����B���z8vg��6�>xQ.�T�������L6]pS���v~��g��T�e�byr����ϱl���n6���^T��~O_�Jr�y�^V��6�Y{G^s�,����u�f�)��mf��"��^,|������8 D�@C�����\�7t$������4����1+*.=v��8v�/pb�Z	<