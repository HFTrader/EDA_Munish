XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A��.�ApC�p�$�/Z|��(�.�Fn��o���;�s�9W�b�/�K>-|��O;���Z'�m��No0��:���=ײ�d�w-�ak+�	�%|�k7×�w�s��+��<r(+8�����g���g�r��g-��|�0*��`�\/��n �}�>;��~8m�o:>\A��4J�����֧2����ձ�2��ȁV�����G�	���&���Yh˽��OL��!HV�k�r�ס����p���ʂ0H��i�ss�Kw9���pp�9��éH���l�~�%<�ǟ��BS#}\����!}i�?�fQfF@c#�bj)[cS�9�=�ILiۘ_�$��F�[��Z�JI�/{�\.�09�&�:�xD;3�oF�Sm����Sm�r�;��o��m��"I$�b���j����������ߟ��z�m[�a���o>�;OJR�c���Jc'��w��L���ڲ^�Dsq9�j�G��2���B���#�/&�� f10��-,R_$��� 9,����w�;krr��Ѳ{�[E�!r������i�7"���F�v���p���|-�R�|L'O�&T±��֭^9��<������V�3���=��epM��|n�Մ؏�T��#P�!j��7#d�ޖGn8N�/�Ϫ�W0f��Oه`���3C�\N2y�Se��""���C��>6Q������X��Hs�t%��= 5]?�]��O�Mp��ex��e�~�R�����MʟA�VO��K;��]��XlxVHYEB    17c1     810J�����q�-�9�����7�_J[ߦ�%M��~�ۦ���%�������z"�.�c���Wk�<x�Er���fw��_x�^!Ѭ{8ؐ|��d�|�[�'L��L��pdh.�.��w8(?� hXn8Z�պ�GK4c̓�/������<��L���
`��DA;���d��[?*y?-j1�;)S���> Xk~�^�%M]AsC�-�p\�٫'4?ܵ�UѶ��G=_��d�5�@��V|��T_h�q�^����9q�yAV�S
����-������'�����J��O�~��<�>�&�AW;��@�2d��V-�P�FН:Em��'�P�G5�%	﷭,^��J ��e}*����\���ڞ��h�,"���9�.�
oJe``�>s��)���}��G@��M4��4����V2�a�2zd<b���Hd���%��(ݵ$���ŷZ������`R��!˩ �`9�{0l���Ć���y��Э���';�RJD~
�^�,Kbai��/RT�7���̀D�G�����o�B�FFA�CqA?�w�e��<��=8�ߟ���:o��N
�G��m&�C�~(9nn��6�yiL�)ĐR�]���4����A��QE����A�xI#�T�s��ت����p����~Jb���
���ϱ��cA�p��u�
��e6��aG;�!��.[�e�/�E�?�Ż��\��8�5�)�B���B��ЊL/)mWȃ�I��š[,:!���^:Щ�����%��1K��s9|de�B?=�����4j$�>�IT ��#��5�#�,�C�J5�䇝�m��"�
�}��;��7H�2��G�t�X H����w6�-�	�[�s���'Ug-!"X�t���w��XJ�ؑP��0E)��W��9SS�������g�0�D��c� /�TCu`X߯(@�?J��K��x�FJɉ�У �]l�l��A��K�a�����(x��-�M	����ԥ�԰Em�v,� �V��\�Z������Mx2^��
���`5.A�i���pw�� BDm�o�y���1,js�v�~���9���!�Xu��9bN'�P��"�8g_��I��>��D�j�<�.��M�HVu��~�G?��g�*�7:??���Ӊ�)T"��_��W���3�9�j��dP(~ʒ �=��-vMj(M��b�h�zjT}�����&ʥ:s��"��4;?@#p���I�뮮�4��frD���h|gi� F��҆�9��(��Ҕ���¤|��e��FX�ă�K�7�Mn�N��'l �~��1Ru�T��7[#U���O�h|*����T���AG���ɂ�=L�d�ӌR{L�ײJ��KM�IӁ���=�d�DߖM#5�fę���"uP��|sR�HMqj=A*���	���{�w�1�7X���i
4��_��V�U3j�O0�`҇`Z6�X��D�Ƌ�"��&���hQɰ�m���?�I�lO��;�\U��Ǜ̽�p�	��9���a�'���~%�Okȉz��O*�#k�;�;�~����jB<�_��܉S�G0���1�0�j=Y���E�r �$|��_JT4���_���������giv0��Ʋ��tm�P.���D趴3ԡ���A�-�RC4�ʅ��ֆ��N���VkF�����Ҍ��3���}�d��W#m`np-��S�п%kJ��Ӆ/��"^U��lo;;���=��O���|�<���I8�����<���;Di�9Gi���9ڗ�q�������U�9h��r�~#��c��XJ�2�5.?j�;�ͨ�urcT{��P]��O�6G��RV��5UB���x�I��ՄB0&��8V�i�]ZG_�i�O� �e�p^Ɣ�M�+9A����pH�,���]��wC:�O�� ��EyӇe���a'P
<��i`i�!������~,�[%���AW�Y`��Ɔ��Lhkjr�kZ��&���E�q6\�$g�/��ǻh���aާ9��.觌�ȗ�^��t>(N#�ʁ