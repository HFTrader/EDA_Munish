XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'\�Sur����*��P��5t�bU#�Y;�`G�4.�	�ߘgR+��K8���u�U�q�yv܎����X���+�f݀�eW��*\�Q��W����-��\�ŚR�g�7@����xw�O��pU]G��}�>ZR ��vЏE�~�2"xR�<��=o�Z0�^z�@�(}K5f��0�\�醫��٤��?L���;н�>�#]���g >�ѭ��`_Dbi���rKx[ꯂ���B�{�5U���^�y9 Y��V`�D溥�������&� 8��y��-��	����v���T6�қ�I�i��m5-�W��e5�W�۵!8�E���
�i�/����)��Jz��{3��xLf�c�0��:�)���Z&��AME�*������*Aݹ��\��aU?[־���|O�ˌ�`;�n�������U�Cr�;��s������4j�͘�79�V�C�k���?`�'~"j�L�N�������לOai����zf"!\�ޡ�8간8�Cn��������"w��Ïi����g(nlօ/#�96)>�0�a�T��p]n�܏��uY����i�$�%.>T����f'�r�1.1,�5F�V_v?z�#FR/֮�a郼�	}������;���bX�m�ƶγ��L�xK6r��2u�P�Bα���D �>��s�?A�ŵ��s_��!�Aê�+�',4�	�FjT_��bKb I�^�*t1@u=���PsV�O����2�,j���e��-�%d���b�6XlxVHYEB    17d8     890�s a:�`]In��fQJ$i%k�����͐"�	[���>�E�IB>L�k�,�貞Q��k�0��r�c��nI*���2ҩ���q������E�Pc��@D�'�F�|W0�caO�0��U<̵U��-bx�wzZ�.6ȚY�l�c�Q�n��']z������?���9r&��F���N�����
t�G8���m��j�٣�>�~�㩕�\��y���<>[]d"�=�D5�D�����%sV$�g���~�#���'E�K]�.s�bq`P����$�;�?M���<gu#�8"�\��ys�QM܁�f���-�|O\3�
�8��s���VI�ujIB|�G!A��ͯ��8��C��� ���`�f��=|�w��k�\�2:8�$���㫊oT�PB�O�K��pb��b���_�9 �]y�����ᾝ)�I㗜����26+�|y8�2S%b��
Y\�D+�a�QdE�H��'��޲����C#��I
z�Ǐzg�07�k&�]�DrxZ��J��&M>9t�l��D��s+Q=D``�OM��c-�a��҇�3}�}U�O�(�H"g$��É��[4�l	��,B�?������k!���pl�;b�į��r>,E��e����U� �A�b���GDoô]�tJ���:��Bq�B��2�(oy�$���s�I%2\	]�.���$S��U�d�zQUI�	{��G���a~xb��3ܣ�T杕�% ;e̗�)����}�]JO�и�ዕG޶�M�-�]�"Qh�Q��� �C�����S�J3!S��z����%o�(�����WFMЎ��^َ�?-ݥON�w�J_�vVO���1M 7>t4�j\�K˅�e�3s���!6�EiB��g+�x�&�@e����v.}SR5D��l���4���Ĕ��Hh&Е*⭄5X<�@��IMX��$d�gL6�=m�b?#M$P�|��ɟ"��D�_�4��ƿ��F,�[�oS���Q#ؚ���K���7E*�Dƅ�����ᦤ�|&4�����I�ɬt�G �~e�o�m7���C58ѹ�Q�Ζ��\*Ɠ��0v{%S��f�&���ʒ�GB� ��:ڕ���NFu=k2ӧ*&�%�04�>�?�Q���$�R2�D�d�|c��"������4��@u�+􏱖'�q���Df���I[G�V�`F*Gs~Nh+�ŉ��:1�r8I��!J���I�F�|�o�)�Uq�y�@���<��n(���0��F��:�h%ѹJ���s%�"���U��mug:�-x�\�����[�m����j�\nv�A���s�	�[��`���H�*�ƷV���T<5A�D��ވp6��m���� ��]��m���tW�5�����r�8
�uz\$�<7�L:��l��'�zt�ʔ^[}�=5��rh)�-܋D�}]֢T�yP��Sڱ�5����EpU�Ov��~ZzF��p�o�����^.wg�>��ab�+	X�ڠ�/cb"���%���LͅZ<��	� 6�'��r��͒Q�% 8(Tm
^F�����YY����}�E��C��t����V�{�Xj���]T�@�&V�8�n�R&���M�_ ��E��Ŧ�E"���߆jYh�T� �D�� Lk�bϪ��eKG��=��Z�]<B��RXYi�jҖmL��))�}q?�̛ևpDi�+�!�'��N ���@�6ǼMU�t�P��d�JK�َ�Zt\��|Ѯ��T�ͯ�����mja�}�ӟ�F¶��R�Jh��=H"�A�|)�Ǧ 	�b=&\��*��H2&���m� �'��t���n��K~&=���g��4>�����醺�M5�i6��6����n)�f��{����A"����J�6HD���a�s?��]��n� `�0h�8�P{6��|�a�dlʃ��?��,3˴hx�H(j߳�]y�B�T�Fz��q�+S��3y9*7����:OK�\��r+z*Y�&I���f~���̜_�&�<+	�)E�G&MU���" {n���	I��ԍ��k4����B_[��~�2`��F{ȁ�x�[g<y��޹"�-����b&��Ǟ�+��F���zTbN:��&�]��Np��P�&�$���`����[���	�o!݁G������U&���d'