XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\��%�r��50�D� F<�^ʭY4����ļ���@�������lXmW��SѬ��J�q�\%�����ìI��M�C̈�4^�5C�'#��6�N�s���C���=n`,6GHܧ���@*�f�a���L��d��E� ���]�0���[��j�CHi?��'T""�x���Ĺ�y+r%�w*� zD6~U{��v��������{�e-P|~u�|����Α9Vgz��9��թj�5N�i�XP�����E�Щ�9]�r�ER��FKɊs��B"l�.�l\�C�5�0�?�N2��ݴ�B-b^u5�ȡJ4� ��.�8^��N%����u�#�tq~亱�����Y��N.��F�\����O98ʁ{
X�e�Ł����`i�~>,��3� �#��XWY���}�7����R͛뤟M���~�{��^�N9����#6S�zP]T�Nxi�
l��6�Vz$���;c���k!��ET^�Eb�q�'%�_&��������0el���i����#/ǻ� M ��*�)�	i����aB��U��wT2N�A�����²���Ϭ#����G����3�⏡eL�{_���/�k�͌k�k�)�Yυ��j��^����Br#0ĳ�4�j�\�z:C���\�R!�� A
����C�0w��pH1�o٭�� �$��n������13!�5���������sѪ�	a��=\�.��m�{m�����i\0��m)�=?�J!����XlxVHYEB    125b     750�K{��=�K�"@��|��p_$�������N��k,i-���FE�B[�3��8�'���*k���*�j&��ơ�LJ9�d랛�1��n����L݆�[ E�ng����Bs�L�E�63�8�y��k��0>Q.��^��­I��U�t�H�!y���^�\�_��Q(�m�脺���S�Z�_�1���3��]�vsu�L���x�1�1\������8��:��'�}B���-p?x@P����\�3�am�o�mv0�7�I&������>@L��4+���3���P(_��������lG�/ujPjYH)e�h�Ď�L�	�A�U��(����&X�'+;�WX �!wT\=G� 0i�Kɀo��ͣ�V������]�`�L�l�f��jJ&Yy���#�wV�6�sƍ�S�5A=�Oi�V`����_bC�d��q���G�*pRn�;=�!(��q��D�6���7�|zB䦽Vy����%�}��e�큊�:?����W_XG�����x�!��h�3`v:1�)�{�j���{��[!�ZuS�醳�q�9�^���&D�	��ơYG���W���L�lnL��5V�������\F�u�5]�VM�!Pk����=?�d?;��wa;"������]��)\gǍ6]J̑ ��;��t���h��v1�B���G��}P���T���NK٦��G��`"�� �d�쌮�]ΐ�����cE���:T��|
yȖ�N���/3=*G2�A��Y<J%������)�71��>�v�j��X)+[n�:M٭s����L>��"�u��"Q̇cn��4,�e�y�ZK�~	޳��B#����Am0Bo��,�~��\y!��88�.�L^a~�a%�	��-�R��,ߟ/8���?�q�AoG�y�XX,�c���du�8����(�7]S�V��r��nѳ���bp�����ؖ��Nx�15��I�Cw�yT���!�t��u�fD""6nG4�۹X���2��X~hIW؉��<{��嶑�J>�w�@\~]�"�D0�0���q�;߉k�1���LYW��A=�|�O��xR��Ģ$�hw�h�,�b��%���nd�Q��\u���W���7=x�ʬ��.�Lf�Ӯ<`���1�O��?_�-D�-��2�Z{.���1wQ�Dʨ�bn��m��/a����S��H�	f֦���Ɲw�%���+L>��#_#�pL������c}lo[��[}��/g!JP�z瓭IV�ސfVI(4��%�)2j���b-�KW�v�`l���\���C;�x��Lp��(g�f^�������D�1����|GT#R@�Z&L��"�P0�S�@�;_a���[Emb������]x7�˲�7�\׻.�x�!��@��� J�X���aZ�Jj?;(���M�����~�}j3� H�����@'-쮐&��x��}�[+�7���:�n]�]ޥ� kiv�e�2�{�ߡ�'���-��ѯ�U��QE�_��-�NÂ�{�B���Z:a(�;b�`�i|��j/�Iؚ�8z���<h��b\m8;��n1�ĢW�)���a?q��o�����0!��"��w«�aZpv�C��s���%�Aչ{#�GU�2������� ϴ�ް��,�����g��_h�����P5|�@�tg���~\rr;�M��2�?��GD��{�0�Y�܂�����aĒe��&��t))
�/R����u�]����X��3����gr��q�k�Qx�g!H�J��s�u,�)�V+s	�'���-�KCP��6v�g@����>�@4��9�>���[��[���$�_
E���cX�