XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���tD���:������c�u<9
��x�=EԊ��#v����#&#�^褒���<9!$��`�+�(�a�TU'���rWV����nv�ż&"���_�f��ݤ���K��0Y�i��z8���l ��@�\?�<�M�ع�H�-p�A��gP�M������e��*�d�+/�49�@�@���x�1�NZ"٨�(sվ�3�ނM+N�NO\Ӛz��u��a{�!�����(:Xx�D�ǃuLe��)h�6u�k3HS5%����������Iym�в
�<��4p�ȱL&���w���Om�nj�%9㹮�L1��LE��f��YZH�}��P9'#|	�#��[F�b9�Yz�TA�T)��
z�3�e�J�b�����g$����Fqi��I_yuĲ����p'���N�X*���}��cr����=�=�)����)ox�S��7!�E�\�7�a�������g�Wp���Ϝ-���Cb�[~|�Ô�!e}�3��4%	�t�b���l�	������O*�g����@��6z��0gD8e�v��^@$����6��!⏶�BUu#�E�<H��)��t�SY�	a��� &�U�Y�o�J��?�KgY9���2	�.�H����O���.V4��
^6WŁ`����
\�ZwK�١�����q������_�b�w��Y���1���[�Qę���d�(������wA-jLt*�]A�{t���N2"��ov?�dOC�)��V ���%�HXlxVHYEB    32e2     b60�3l�҄����]�8��'���,����1��Vӟ�jy��g!�E�F�g��L��VҵG펄4}�5&ř�!(�������D7\;��Tъ�w=>�o�h�s�&�U�A(2p�a>��_�M��J2��1�(
�'��,ԢG+��h���J&�إ8�B��6T�r�ЈO�f\���N�7-=�1B��P7}F���ѡ�D�+#�n����`���m��T�[���$��%N@%��#�ۘ]�/ԥB|��r=����7<'�V� 5˞22�&�W^M�~�Ҭ�C��)�s݀ ��7��!��@�_M�}���q�M@��ys�Di�6*�h4�����Bq�������t]���k�o��l�zZ�#i+���1�v����(��	ҕ�h��o��������X��	YǷ��� ��d+��{j,� &�an$���W�ȧQ��B��{m�T��Ȝk6R�Px� ^��+ �y�g�2?!\��c1���3��h�I~�Q�R�U[*��8y��3q��D�wL\r�F�����='*S�L���)�WK�)8�������gQ{K��'���o[0p�~���p�F�>]�D"ݿkrr4��aQ�����$�N�h�_[�!3��=Dgo+���U�%���e���ɞ� �U�Y���I\5�C�����pkԞ�-a�v��*�iG��ci���!\�_Zu��Q�+S(h��Z���Ĕ��[*��֡��yV��h�2��A�~�O](9/�^��v�7�����,�֔�� #%P9��| ���O��V	��ߊU����~G�Np�u���@g�0kHTF�%���I�����v�$�$���UX�Ns��k��\[��w���������'�����LS����y�{�b���p��X%�����Æ�5�i{K�:<���]�U�r���Ga����,�@��I��{�<������:Il8m���Z����Wٴ�ƈs�X"��7�oC�$0ת���3�UPryIԤ�2#Q�6�HU������'��݄)����#�gю-���YC��'�C�ޥ�@��^u��sd�9j��K@�4�U�Q�Z�@!�d�?'��@o�.�!fR{��W����[j{�/%��<���$ڦ3Q�?�������>��_)���C��U|J�Ȑ[�=[��+ �V��9��`�B��2�����<�܎�[P�tQ��P���A����g�sW�.����ረ���5r�w���Ow6�����и|X]����-@�ې,��1�I�E�C5Vm��< �oN��3�2j��T�޺Fʳ�Li�F�O>�ؾ6'R���7�i$�2��>_#j����*C��\r�A��^�ۿ�O8c���^r�?��pwC�nG�s9��
\�d��BDb�:(A�i��{@��;���[h~шK�l�߷'ͺ�)b���બ@u�-��+*�U��(X 	w߳X�e�ٹ�e]��<�?�px�3#�ᗘ�l�O]
Y��c$�	�N��{���h�d�؏}YE��b�G�{,8n�k�Ƒ�r1�%��%�{n��!��@��>�z���e	�@�!L�3`le�u�̠ռ���q���������Sɪ�t�_�m5Ǡԟ&�)&,KO�����PO�^|�~$�D��Q�*��F���u��o�;���v@�d��xZԕ�ک�O)�I�
����AEK}�-�r�M���Q��b�9�HV���rga;!'*u����4BG;X����7E�0(�������1?MR_j�Ң��6zq��r�V�k�*���%�cOM}]�����monv���_*�.��a�����_���8�O�ӌa�n֐/#��y��J%v�������xM��Ŝ�*UЂ���F��M>!��#�N �K�5Nά�g��n=� ����H�m;��+|P�n�z��X��J�q�,�S�<m�Sc8}+A9�[�ߧ����%��cŕ��"�B TQL�H"R�n��<XY���Q�p�o��u�������G�����
iϏ�z���᭯sO��`�'�['.�eT|� ���ul,y'$���}�{,u~����׊��x�Z݆���-;��N���2�M�gh|�]]�'��-���Ԋ4B��3V��C�(�ܘ���*���H	yP�W祯�R{�C�s��K	}�j ��a����O��Q��5�n^b{��;��g�Y�j��n�ȉO��*K��Ž��	v�����k.��G� �{�0r�����&;AE�:��|�D�ye0�{��J!�&ks5��)�(��у�D!��f�7�"u�v�N��*X�Gε޸,[���/m���㰔V��UK�t9����;5i��?��m�-��Z�,���IV%�N�~�.Y��5d@���8cG��A�~j@���"�)��S�
��CWsZ�8���Q��\j��7`d�-6)���g��ۨ�b�`)i,H�6�9oI�}E1����[��\�ؔR
X%�g@
��Pʔ*�Ic�,
�
��W�r�F��xVӎ���7����ĵ@pu��M�\�
����I�g�����b��pnQ��te����cb����W �Z:GB��H�-�g{=��|���*���:��&���R�1��w>�Q"�*eOm��.�_ʆ����N�i~26���i���܂>�s&��8sIܧ;�ı�$�*1Z"��u�Ǒ��˳`�M�K�>����"� �$ط�w��B�f�{���1�O��ׅ(5(�'-�?����h� �
5�晽����RDK�(A7}x	G� � 	����q�Z��F�^�+be>�X0�퓎��a\pp..��̖ζ����Ȍ���