XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i1����f3�U�Q��EH���Sn8��/�ߞ˛�	�_�B��5I)"��'��*�G��V�S;�������[LcB`=�h� +���Y�0��m���/��9AR ٶ5B=���'�i����c̲���&��h��m���^>�㞩�@��؜�~�][����S�}��.���B�J2>��L	g���j�]��,�ARD���. Ҷ��a�2�-Ȱ��}ׅw������kJ.t��SNg�Ϟ��l ƙ���j�����4��A�lÈ��"W�#!ac;�Bd����Mul�Ǉ��F}����� p�
����+|����5����5�5�{��O+�fD!?XWSfc�=��L�lǫLH���_�>���`|;(�_I��^�!��ٵ'��b����q�ٽ$��e�9_�tvO�@D��ܴ�]D7GܬT��͛8��s��wTk�T��(�\��/j��L�_@���D��~�y���`��T9Ѣ�]���e����>�]��P�i�7ẕ�W��%���N"�h(b���+�4`
)��#J�n{�}���&/�V�_}�>ሕ�lJ���p��l��T!{��%J� M�3IB�S�X
V�ǽ�vE�1w<-H!�J�\���![!��Й�É$�w�k(�v��M���Dn���.c��T�o���<W_b�4�	Y��	�Jq��k֖)���.0M��p�(=vU� �([h|y.;��Ж�=���g��`]�v��I��#XlxVHYEB    dd8f    2160x���$�3Yd?�ף�]���ւ]��Q�"U@�5��!V�>U�|��dw�������1��1��L��F���fVSi��m����8�~"k?fidZ�.FS�����7��aԒ�O��K-j-#�tM�ވL�ѡ�tl�e�-�M�=h���k�_����F�yA�G���܌Q<�+rb���$=E��)��bq�����zЁ�?��0��3�%�B�wéb��ZC�91�Q�ܼ�o�l�9���U@+�y��pù��d*48SZ�&��;2ل�)����i�cnt�tݎr����13�����Ĵx?eaH�Ax�I���>&�e��Z��]M����:�}��>�4?ȿP�u��ґw�tg����J)���EŃ�Қ��{X!����fos�΂SˠH�	1�n�V�y�:=^g����0�%Q��C��K�,]oC@�A�Xj�����t��`�d���]���6�qFS���	�rZu���x����,g�����[AG�j�x\���?�g+f�UzP{��<W��$e�3�=�"�)l	!%�w�w";��IҞF����
���*��}��9�B��������wpD�I	0��n��v=ڿ���s�d]_um����y��d��o�S�x�N(�{��{�I�ʷ��ɩ�mu�sB�V'�#1�z6#?h�\���|aE��g�Mx��;%�4�D+~t�8�����L�\�Zm������E�wA�`�A�z�N�xت�½0�b43BƳ˾������C?����2E�D���z�V�$�TC �ټ��D�"���@��i���Ct�Ɲ�%���F��k�m5|YJ�m��2J��o۬h�s荠��3�G_.��Y���.Q@ʋ��N4ڪ�1�gC��#O��
������1��<c��CΟ���F�s>kB�ƄO�w�w530"���X�G̾4��<���5��[h�z���@�	�����Y6�X���1b)>n�#CS1�l�V��y��"�i�󞽺�����W\�`�ę��#^����3�W�EM�L��%;�U�{���S���v�T�9��x���~L��jB����`N��R���ˮO�I�`�7�7 fWy1:G�J�l���<�,� M�Օ���}��D��ύ�B�)�Ap����1��
Xݢ9q���V��[n�;�J7�Q�4��@�)D�s��_����u_aj��`��Q̉?��6FuLv�U!��Ӡ�~P륈չ	`�l.����G�^��*����T�A����F�GϋFo<��À�񈰨J,��Ú=m��oy {Hl��w1��<����~.W�6�ۗ{���"❞�H�1=U��f�G��{������ݾ��T ���bm� ��'h6�������Z	>� "){iw$̤�>K�W������Q5έ�z���ה`g�n��e���k]U]x�]�����;�����1r�v('��E�^�%�e���>���4\dx�2��ʢ	#�ƘWv��c�#������L���F?����Z"����\"���0s�˜a�M�_N�$h��|=0�+r���d��Ű�j�����x��Zi#4C>-�r�]2�[�q�%Mf�D��Υ܉�kl��<�nWV��Cy���]��B�a���C@A3�'ԁ��Ek6�H44J�dD㎾��fk��m%����="����HlvY�lP��f�D;�z��Vl�fX�;������bM�+A�W�,� ��\V�5/,�#��_�v�b�Af��������~�+Mi�h���͘����K\��Г���u�6����]d�eR��a�:����:��1�o6l2 C��[��=v������������Xv��oc�9+)�d���W�h����"�۟l�4;��-6_��qk��V��^�KQ���P�&E�-���kv��j�Z!Yi�%��[�WW~1�k�ǂ=��cN7�$�.��F���r�����W����efБ��Y�3+�׭I��_�q2ʣ0V���\���g'�>��ʽ6�Vێ�5�K�RTyJ��:�o��1��lm������2�����H2H~A���Z�^�;;�I3i> ��O�����O��Ō���1���JM��7����D���T�]xy��>JNY�C-�Nٽ�+|�IT�#(�i��^k�w&	�M�DI����+���(+�}͉\MeZ��e��8��+-v,��
�Hԭd�E][F��loV*�h��n�z>�MF��fC%�6�3҈Ն����<F�Μ�S�ըD��`d��П�"�O�ef��g� l=8o��%����Ld�O�]����g�k���4[����4:PR�}��j��5�v���,�l"�r�KCfg�?�ģ��?ۈ�w�B�ކ��E@:���l�E_���!"��KG���h�,�?*u3�ӌ�@ko������ �%-8�����L�������!$x��dX�V�}�M�P�ӎ�է0,�]
5g��P��I�p3��k�=��K�	%-�^�1t[�t��X{�[ ^C����'lF�+_��<�-EK��v��k4��Ӛ�|gb�<c�b������(G g��u�y+Q~u�kd��,�6;Β�rf�=4O�:/��M�.�e�8J3��Y���Y ���pZ��R]p!J�Kut�H�����d7C~R����R6`�{|��S ����h[R3�p�D"��5�%�L,���@m���u|��NX,^�]���N}�3۴�븞���󯧱�.������{6�&��-�r[9���%d�5�@9�-=P6�2wF��؜཭/��Wz�0�dYW��r|�v�{���k��a}լ!3T]	@E��7�,�t���d8L�j2Д�u��V�1>T���[�0P�'��/�ˠ�C��	I�r����ah�r���f@S�#6,f,�*�F���
$���EsP���
'YB�7�⏋�Sx>^�[mS���~� nc��px��X�\0�,q�[��Iz�&�����f�<[3��~ �/�4y��@o�Z����<*�h��֖�/�K�
z.3��Qrq�u��k�Sr=�iUs���*��9%�7C2�+�F׃�;fb�<���ʇ9�{2���d�9w�5�q#�#���ܣeFu�d�/MΫXK`{����s�����7�E��gTc>��7�4�xb^���=��s��� �r�ANI�,��^����h�m��%�K���ބ���|��o&�N��Z!�������L����]ǢV�*z�RC�X[�0�#�Vw9UxI�>vq�t�Yi�#WV����,3U�PNȳ�8��!�ڮ/�>��<$k���{
0�A J$]�����te�~�o*�7UQE�!��粭f1�5���]t
\������;�CG	�K��z��תv��w����-��I��/r </t��|��N����ݓ��a+R��[�
��\t��^�3��úN�=�Lv
P)�ϣ��8��.e�r�y��?�Q]������mNcR��ǭ�/:��s�^����MHݽ*቉t���D�#p��a�kKW�WwvxJ������x�+2��H3�duk�<�N�x�W���]����UWl	E&�}��c��t���a���;��&
VdC�M�\:�y���k��8Q!0.�K�]o��KVj��MD��}�}��^��U�������|w�/�2�ט��œ6��L`:���<4��N�s���i��"�c�:]ɿr[���Jd����N�e	�{��˵�s���4	뮥q��Q��Dc���e��bK��wSS����s"itj!�/Gv�	�VD[2�D`�z���JM�X�~uEg��`�w��jPQPbLe,�d�ф��hĵ�<�]�%�T;��IwN�rn�ӄ�˜c5�Қ��*�*����"a���*��s�an���<���Y��B!������3n��;��6�R�̐���.3�K�c�Y$�ƇOw��C9�Zcx�h��5�Q��7���E����	H�t�|��w�y�@�@����Up��X
C��䫶�*���xt5�-�JE�������bR����;w��w9x�}�� ڀ��5J/|�δJ.�5�d����N���$��x��Pi��@�k�hȢ_�����}KJ�$L<��C���"�$��.�\��4����f��>�j�1��_t3`;<�	F��uA^$3��%��;���[�-gӲ�JeHo�Z�TeF�\���q0ۃ�d�jCqH2:��O��'���|)cۀ����E-Uq{g�&	��M��Y0��~���45��ekv��$�:�B�@����J���UËC��.��o��ۆ�'?�5��[�0i�`��֧竗�s�^�yKC�!(G��w����x�|q�	<����ZJ%�����;��@�I�;��y��\ �VW�Qޜ��ڞ|�� $���Q�s���RrX�ik�ۼ��Ã����v�?���ܓ%�r��d��db=F^k1�d"@uG�؟��4LƮG��O��g>�f�pI�0Ky@8�OGQ���.g�n:�/V�ƬE,��X�r5�D�2t3Ɲ3�!y���2Njr݄�E'������A�CPm�����2u���3��bY��-��������z���p|�5�a��Ґ���
���`�h�(���O|\WY=���؞D�����h�>��-�Bڛ�����4�}�ÉP�����Qc�y��'��0�z����Z��� ���?�D P:��Q	��
�t�s`^h����)+�
��{��?uO��yc�"(4�_�E�LN�T�ƯyP�9�Ht ��~'!A����W��X��?.��R���*�m��9��8�8����$����|B��@��~n��X��J_=�`�@ȑu=���%c�/OQ��إ��#KE�������7����ֶ�F������@�QL)�q�MfE�Nþ�?�e�N3�o|�[9��Ȑ����=���煄���Kc����h�����}0�Q*3/ioT"B���!��!���3Ŋ���9�P>�ebd�)4�07 ���n�'w@R�Y��{v"�ꢲ2~A]i��~�UMpq�0���d�B�!�z�C��B!�+�x��N֮D�;X�v����]������n����d�sCp�o.h"8zCއ�%���^f-�V�_�1�kvˑeX�Y��i�l4�¦����1L����Gl�p_�ZMy�d4A�0"B�x;+7٩��Y�әJ6]�X9����J�h�T��P�J0�#AZ�i�5%����GT%��^��^���>�)޲�jb���뿭��q��!��w[�\�qY�2.$�F��0Z��A꫉шE���b�߳Z���+���`KY�ӍW�z�#�M^-%�������O���� �X@�@&���)��u��OX^����r��O6q��ݳw�7O!��
@����a/��1)� ҇�ul舓`����ʉX��vbR	r�����d�u� ���̍�d�{�87e���^*v	Ov���*�e��M�[���P���7x���qv��6KR��4��߲��N�p��n�%y��ݙ�;W)u�\0��f̩LO�����6R
��͂�i.�l�GX�����u��0��Oc����n�uw�l(��9j7+^�K������?�.�ҡ3O���,�2��R*��w�]Hq��7���r�o-A���O�@��Sǈ�b����!��j;��/�����MYtN�)AbW�Tg���0,��2�� UF�#���%@~����3�$A��53��Zn���=@~���({(�ϖR
Q��dZ/A��T���)���l 7�`3���΄t����Z��-XLP*��n__c9�`�z�+G*�Wi>�K�m������LF�\���sǒ(��2��j�`���S�>Ʈ�n��r���|o�h��U� $�c�B><�����	JiK	��[Fx?���M����o/PB~�P�Q�7cn!��T�V�ѭ<�%��̏�>,$����i\5-�>�ᩣ�<�g�:k��G��$�`(�.�!�	�	��7���<i�������H0��T>�(ш����|פ��ۮϨK�i��g�:�MP��UM�5�ս��q��X����a��OqMO�ղ*�m�5�Ja&�jJ��{<�{����S+wm����
��0C�y��h�l��z��l�n2"t7�-���,����[�C�fi��E�Q�U�����d&w�@�F� �7����0�u1$x�R������l�]�|%ąDo{���LG�"����O\�eP�>J<bI���Kp-9�{)��z���~mq�3r�&lܝ␝#Sk��q�����5��S���*��vH?���GO-��+�=ڑ���	xc�gl�>���w*h��|�>��)�:wy���r��)@�V�Z�ȖN%�Y�B���q��X"t ��}r���T�*Anv�P�;]����f��,��;y�L�qLs\���ȋ�PR��⌴WO)W�:�.1y�]�]��Q>Ϋ ���,���r��w�ܚ����ԇ����8R ~=:����1���R�5'��{�hd�p��Ǹvo�S,�T~-l�[�g��4�c� G����tJ���%C�홮(S�qycB��.z-o�]]�̇���?�%��IQm�\;F�ԭ:�S��vY"���������������X��'#Y��.#X�B!F���tI�Q�?Y8�-<�L?�X
Zx�]�Bݮ[Y�+Խ��E�[A� `t�^��ڋv;9�n��jQ'��~�sQ4)����� �����k%��,�k�Uzn�N�_K�Ύ�U��<�W N�/��gPH�Ϫ�.���n��-�~�7�����~m~�ۤ n)#�eBJE �`�����!I����@O����wA�"�.��Me��!� :�˫v(Hꋁ}8�3/����RB�\���!MÇ�j�����W�.��=
�$-fL�\8~ֿflz�d�� ��;
��*��c[َk�t��8��Ԝ�K�H�L�a:��ïNz9�W&?��|H(���y�K啱�z鑥Ũ�K;3�#Z%p�:�������m�D�ڬ�����|N(��}�����YS�ғ(�&���G�z��.a1��	=//vB9����*�u�4�����$�|��I��Ϋ���dUA;� *Rp��5�埣)%B:+��ἤ�t���BI�e�xb�=���e\pxGx8���(�$���'Փv"�-iC3յ��u%޿i�����ȯ�̷�6��^���� L��H+��������<L�����L	��!#@�3!�$�Ȝtm�,Gd��mW>�M=�**�v7C��]WR��xx�M%���4�`���o9��谙c�ڲ��� �����n�+�0
j�9)�U�MJ���X	��{x�mߵK-��3��hzկ_<��6���>�aл��z}��=.[����ꗨ]o���6{o,l�gU>�����ʾ��u�y�;��Cֽ����8<�V
���E)3_���qL��m\�����_�&h���/(�2h|���;�}i$��J��)'ѣ�1B��By���&�r��=/�� Gg �3�?Mq��A|��Rjm��k�旅7�D��V����Z
��Y�W��xk��q�ĉ�ͦV�������L����NM�(QW�s�mŰy�_D�.����`Y$�=��%F#�l/�+u��o���A�P�B���m���fs
����
I�cF+`O�9����������ˋH��[��uFXS��,���U�g
eA�lӢP;3��5׉[�D�𻗥�by�7��m��R��B��4�}����=�E�B���۔�>M���xX�S�����\<j�!M&�=Q�R�f�RR��Т�ԧS�I�U�AT}P&�Jj���%!�1~�[B���#���fQ��w�
\��?%��wr�a-�C�Ȧգ^��d3�D�"��XW�]_J$�G�s�ش�����;���f�B���dv��$")��_�n��3f�I�2+x��r� &���ع���N!#�?�	p��|ՅxF*����
�'N��vb��^�7�)������T�#���b�Gm�5��QaD�h�������_3��E�`�T��0��ʏ�i�({�չx��9���wfw�p.|Q���J-�h	������F��}�n�yv�R�Ig�r��y�.�{�oC~ߐw����n�Bp�ӑ�41�,�ٍ�M���s������xo��6B�SukM4.vԳ�5Fv�{��e�H{�&�6�7�m�k�=hBhʐS�<�Kg��̅ډ