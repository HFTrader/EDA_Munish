XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��:����2�SaM���3>��(������ϡ�k�5)�������	�	p�v��ke��|����ο΃q��at#mM�*,d�*V�	36<c�ͻ����Ee^j�������.S�}\}�g��2�ʂ�@���Z6}�l�)dʱF�m�B��TT�bۄ"\"Ȱ*-��_�s��ۃ�7GR���q�[Od!�[s��-,�X������}A���
���������}�7�~�Ұ�"��2��3�Tk\��YЫ�}&F��T�81l	f;9G���%V⾴�nȐaB�h9���1c�EM�8ջ�h�F_M�*w��g����|��ؕ�<�1�~;�툢�S�|擌�4��l��ж�bᏖ�U�Dc4��� �ibl{�8e��$)Mv�f��:��Tp8u�vs����N<j:�����p-���e�j�X�0h�'�=Z �~�X�;�5��e���f,U�Iܸ�ru�fH�Z���s��"�g��(G��"[���3%vD�Ǜ�F�p�K��W��ӗ`#��ͶG�tp������F���!L��p�,�s�i�N�
�i~J�AH�H��t�{�G�͘�r�!��P�H�����n��<I��G��k��F�.��3 ء�����u:�V�u9�Q�n{>3�!�&!���ATlh�0�����{�|ʡ�`���2��~��%�$ˡ.P�D��	��)�B��J�\m�9��d&�>nQ1V,�$��" ��)4� O�/��5�#9h� `$B�H��`N�'b�6uġ��0ѡXlxVHYEB    fa00    1950�1Kg��A�
@�t]�_�L��FR)������Eq���ྪ=7�j�ӻkAn�Xx`_�����2���.�Bɤ�CE?�*�	�8h'�[ĦSN���0>r��W�e���;�L��pZ|�ꞔX�[Xӈ�q�w�.�B 7��@���J����l[&�8�GS��w-(2���8h�&房�4a����Tz�K'�{����Bp��qs�lOVf��Ư�r,�u�	��X�����<)�KV�H�B4�����e��;a0b��T�(�Plçs�B�����J2���[UF����B������4�N��<�u�*�n�D8��S����v ���yh�Y���L���P$����5)���%�+�/��O��I�h�Q����~+�&@,��m�2�?������L���>B�8�|���K"7��k:3��I%��W/�H�-��x����l83�ڻ�d����WO���	�<Ա�&��Qsٴ��4饷�G����Iu�o2�~鍗,��l��
9�'b��\������ϻtҢ+>�tn�PV�$X{��'h���p�W�dKާ'@�1����>Y\�"��A��/ۛ�oY�%��t%�2a)�󜃑WBwY*�%��@�e��:���ޤ����~����i�v~%�K3�Tx�B�9#o]��v��#dA�w�KƤbyp)z�K��ǆ)���H(���6f��u�ȇ&Ԫ^>(\
�G��S�G���6Ct�_ˁ��4a�0����\2Xqc�"�iA�1�b�+�i_����H��{w˸*������	7SI����4��hX��b9B,[H�v5#�QY��<�Q}~����;��k����vnt,}�i�Ԏ�%��w�Q=jչXCs��m5��4�S,�$ɾ����ʁ��;V�s ��Oe5O��!��L�/D���NwHf��X�'5�zUT��
{��[Kr��Ș�����w?�������(� �ɻ'b���Jc�[E���ιJ�\l�틺)7�Tq�m39qt�Dř-m�ä�Rڃ)��
�Y�j����
�iP�`��Ӿ��oz���H����f�o���\�#�)�^��?LG���)ن�T��v��y)=��{񡟃�¤����.� ��r�&h�e$>swE�@h6�&ef���
�ZB�"��u^ˢ6b~;38CdY]um�v��<@�Ԕᙣ��x	�ǻ�R��N�E�%M/1fy (��R���Wym�O��}u�5],�PɵA6��jC���E&y�tO֨Y�C����cFs%0Ѧ��#��!v��=�>cT�C�G?x<ұ���-#m�A���u ����죙��P}I)o�kf{G�kw��C�E�H�Z�m�n�B	�x�~�5P�[�:�_�x��3b(Tg�7Z{3�Q���	y��e�sC5/@gl�Sk�8	��V
w�S� �'�G]�'�A�^���#�z��p�9�y�B��mA��`3�l�<1=UI�#�-hZ=c:��A�˙�
��Y��G��uЂz�z��E"ެ���L)h��qU5���WB�c{[�B	�T��!.g�B)�@%���X�b�b'��s�r�,��4�D��'C�ܶ|�L���j���b b���#�\C��?8~�u����Q��R����@龫�=�Frh���**☀n�̸�v'��u�-�w��|}t�^oUbPۋǩ'H���tsѳ�w����浖�[�J�>��K�3�٢=��X�HM�hSs�� �&�������ͷZ�,�F�[UaC��#I[�ݝ/�(�ض�x�����X���QUd_�F3�n�~�*��jE�e­�Ùo����b�Q�	zF���������'~[]������n5yO�\(˨�S��,A*���N���W�3�zfi.�c�G���`A8!�u9D�B�m��JgNn jaQ��/�D]G���Q}|x�p��e�L���>�X�?�B_�)	��d�pR��K�x�s ����ߧ�L�����Y��7�Om,`Mۿ�.0�h��f����ؠ��ۅ �o0��U3��n}9��#�h�<;i��A��o7��[]���h��|����h��$���%�İ<�=�X�f�P�z>>4��3�"��NP�N��Y#֪��(��3b���m[�ﲧ�Mv���l�v����Ɩ|O��K�\Bo�&d����0$<e#�{�+�?2�%C�M��XI��u��7R�	�`X[+�i���f�P���蠂���UH��ui6}���:f�A�/Z�WMW��B��i���u)1�`ÐM5��]���eJ����mqF��ifjq��l�n�~X��|� �Q�q���>$�:�n�q�/�&�/G��7���G��I�jC�-�@�{�N/^A��J4�y¥P
)Kt�TҮc}}���-	��<��� R����mͮ9�՚Q��9�c�X+��ϊY�3�!ZA�X�?�����"U�\3�X{G�t�UA�N�I#Z@q/���`lcbX�?S<�u���*h����U�@8���Y�)t�z��,9�ů�,A��<v;;��*�(ĵPEc�D��7Iޏ]ќl2,�Dva!3�T}���wg��*6
�+Kd+%6��*�a��i�����p���<A�b_wF �� ��Z
�/�iU{O��-63N��D�A)��7�[���`e[+Os�n��vc��{y�cw�����Cx�A�%�1I��5=��i����e$Di���F�u�A��b ['O@
`��CU랬����ך̷*O������Y�ƪY����I�ۍ�+�+s�d,��I)�{�:�R�yل@�*v�6��#;+��v�)�$�3ף�7�S��<��V��@j^�n ڂiw?���,ϿφXr��@B̭�¸�R\\��>���<�?@���	���(��a����>���K��L��4re_�B���r$��G�F�P��;�v�i4������s����tE��ĭځ��^m,¾č>-�ث�W;c��e���M��|���mUn�XҞ����)[��D7c�?�Lұe�]%�u	�?0��/��T���t�H��1�u8I�?�Q����y���P.�r>��)zp:m����h�����C;ꝍn0R��٩����hgV ��я�`J�ף����|SƯ��|���bϺ1˹Y��Y-�H��%Q=�b�mE�8̼���v8�q$w�Q����h9!�Rb���p
K[T_�2���v���)(�Zǖ��Ȉ\K*p�0uB��븿:���H��V5����xǭ�LĔ�%n��O !s:^ �ԅMU�����@��*��W��� ��ڢ�0���@x��%���^#�$Ui��^ �Q��L.�>�qR�n�5 ��
��=p��n�gd�CJ8G5X���p�^; ��QO�G��s�06tp����9��멖敮ٛN���s�˱��8�a_==ɀq�O� �M���?�_x���/�#?.W~č�l�i4Y�2,�6\�3���r�Me	Q��ֆR"!��3i)�p_�C�IWȓ�gu
�(P�t+8>eˤVv4!Wzt�Rj�&4��q��j}�q�� i����H��x�ï(��U܊Z".��"�g�`���Ӫ_�v��cT�$��G^P�y�`}�P��Px��g�Aj"7�g��e%O�U_��8I�����OKI��5D��C�������Ǣő���A�0:�w��',����	�R���;G@�=�/���'�{�=A�����c8��a��,�����w|U�ї��I��v��� a@w	N^�|u�&)��ǒ���u_f�65Df� �
�z=�7z-��׀���}��^\��:��I2Vt��7$4fXh#E���Ha��A�?�Btk+,6Bv#v�U9N��u����<�Q3�Ӕ�R/wz�h�����[�_�	��h�O�߫ŋ�y�&PņOU�w���+���8x�ڋ��� }�v]��\P��������3�/v�����C�m�w���Z̥���K
~�.��hf���Ns�f���.r�CW�����>�3}@7e#�x6�Ƕ����k~��'�`H��'�� �Ծ��\���D�eU�ej�VKLP���DF ���U>8�g�f��7[�Q������?W�]GS�͔ACLM4Aw�
C}B��(d�є���oi< D �@;�Z�)��w��x*���kO�&�����{�-\�����������Ö��=0퐢�xۍ5��Vh��/�Į�8�&y��� C��
:Zx��[Lg:et�0�>�k���[��$�9v�����I�TVL'��i���=�L:2o"_��O��~�대����r�{'��*j�'f�ds�e�#�����>��T+A����5�p)��!���	%�����2���I�1lh̸��[A�26�YQ�B��H�b�^�f�Z6�H[��t-�{��u�FW+l(�Vx��
m������qx��<<V]:]?����d��F(�_��InW5��aK�BN��m���1=]�m�#��yR�'|Q>����b��NƟ�?�m���vd��NF�p֡ٛ�U�ЃH�3PI�}|���� � ��b\T˯�\Z��l�^���X|�.і�V�θ| ���"S�E�kq�|$�:Q��&�B��<�8;���Vժ���d���̹S�+D�اX�1{7��X$����,���T�7�?�h�lMf�A��ք��rA�n��u�<ɤ6dJ�j�9[k!m؅yv
�*{�g�º�F��V^b�a���o��d�m��U;a��0�3\�k���Z!��7�D�di��c��$���KO�e���O�jI=sz`�h�Z�/�s�5g�M?ã��)�� �`�2��Zl�Źrp�*���3�~.��Z�wS}�|a��\���4��E�e���?���@����(�4l3?"�X=Z@��q�+�3����r�'�j����\V�C�>OtqÕBF��Wۼ�5ٺD{Ļ��'��(�x�g�:�X�����t�u�OTⴛ�/���Tm^`C1�7��7� )���G������ɝ(�5�p"ᅃ���H���X/�l���5��8e�����~7P�1��b�.�s���fWV_$u�X��=7������$X�{��B���j����+�����<����Eo/�)�`���Ԥ�<	A H'�f1�UO�J�Kp���1J���4�����@}��6������U�j�-���AU��)�Y��k��l@P�3�r>���b)=�i�+��qB�?��E�"��!�1��a
ߛ�*>����Gl��3�O�i��B�|kv���6�X�Ń�)��e�O�H���S°jٹ�_T��ק��%�-��Z��_I�ʅ�P��nN�5�%a�J�F7�M4��[�
`�O�u>1�dZ��6��N2�c���#|K}��`���M����9�����v�3Q#��~8�81\�5��7�|�~c7�<�d�*��`'�&g�mᬅ��%���7��Bm��~�,f��WG�>Y_���>���ub5[�J�E�'��r��G����Qc
��`U؟ci��t��*�:'�^y��1�5*zK���r�9��_��F6O��5�U).�+a��|�C�������;kli#���B�V�|c%m�d5"��L]�ia�K�%���*s�+}�DN�^ٳx���+��ݥBVg���؃���_Y�z��A6и�Dμ��LAЋ�ql�4��m3x������V	����	���J���^Nyĉ�3l��q7�/�<	��'톈P�	����A��S3�#
]�m������ӂ�������:ӹv�]C�	���pA7k���w�~w��|?1��D�P?��7��(E�=	��J�s��6���{ʟ_�~v��t�� ���H�n|�������i�6��N��z���~� U�CLr]}aS�r��8.|�C�%��̇i�T_�zj�B��Y� ���l	��S �V��P���$w����h��,R4C@��.s-���Y|�1���F�>]p��	�O�md,�/��r��,����<�6���[�� 7�1���@��4T���;��^�V�y�I�������ZP���:$�?��mp��:�=�%뙌8)�h6?W6?��\Spg���5�pA=o=�3�_E�nx���m��P$y�7�g��R������Jۮ4g��,��N�	p�tB�`����r����2�[�.���v�1��_]����r=�ɂ�2��Ә�y�K^�`Yn�5�`�>L_Lñ�w�w1	3������k64{�$U�����3�gBW
�>e���~�Q k�AU��XlxVHYEB    fa00     700W�ъ�y`� �Ї���6�̀��!���0�!r�P��F��[��(�~��;�]
�
���p'���\���T$ل�<�Js\����mఅ�����X]�v�	�8�>N�?�A�w$A���b"�"d���|�Y�`�4����I�BNԔjB[:Ф�މ��6��(��wt���_���ϝ)�y�D�ܿ�V���Q5'R�3{������i��X�Y���|�/��z��zMӎh�F\�Poma�b���)�ma��1�_�RӬ��>��e��6D�-X�k`t��d��M��Z�]�b�X��RE���j��i鲘�:q���~rJ&;�7ϲ��xs3����箁~W�C8*	}����^:k��ܚ� !ڴ�iv�[5� ���_���SN���q�@�0��0��x$Lo^(l�J;�������v!�V�AI����nk�❳�u����2���|iK��J͎��2n�t�����ȕaK«����A�NXG���� �dǼ���1�	8 2H�s�N�;N�� `���qG<� �h/���(o� 2 g�U�H2Y��<v��(��\� !����С���p�3�hI�0Ӫ�saH�ɅZ�d�ѡ,��S����(��8L�&mq���i�}ߚ���ہ(&���~�:�s�S�t1ra���?��N��!&��GW��Q��J�*Oi+fG�}��:-Ϝ\M�sS�?��΍W�:V��F�ϖ8��$�7]'���H�<�x
m%�P(�`_GF�Vל�-��}	Ư3��W���yeaEi�R�������eMEj��~�gKi�P�SJ��f��� ��x�F$,���V�5I|z��׽�FQ����׈����L5��H�Kg쯔���.X1L��R��?h�	b�Ei�(eD���}��P��УҒ2�ȱ�;6Ca��gp�#I��ަZM�<����dE:�E��1V;E�^�S_���loK�ؗ��ګ��'����sY�s�
I�sK�Z�jz��&�`#���6����6+�<ҋ�$�0T�b�Ͱ������r�/�1(o��i��!´�E�e��aWk~;�;�j~�$�_�7<sE&>�j$��'�L�:��X�k*8�B�n8A:�D�֨�{A��F�P����6���9�����6D�
�O���;����")&~�-��m��+n:����0E��e�kޱ;� ��~��k��ޗ�U�o��V�$��Pe[h+L���FŞp��/GUo�bT��Lx�k7���-���Pר~��%b}�E�)���4��H�ۇ��� c�Cj�!\4�R"�o��nV&.���ӭQ���<2E˪��`�d��t���Ӗ`Ц�C��l e���W++�<��Z���+�(�DQ{{q]g".��0�n M���#�^�� EkZ�-��fA��⑤I�-�������F2���E[9d�������x��1�ߵ1t�#�I����s GcV]�5�k�P9�����bf�����vu����W5J,Q'��RLXF6�����ܢ᠔ޒ� �c-������	�����\;�� ��[��GE���ʶLu�rP�6��m��B���$����d]P�%�K�9��)X[}�K��}��}�r;4�'�JF�S��m��@R�`�<$�4��F�����֝!��Ք���1��G��o7c�n߭�Y	��75ӿ�qo���{1�l.�*���Y��^�"KW6��f�si�ސ�M��^��2S6�%R�����"P�	.�!򿴠$�Nj��6�XlxVHYEB    77da     a60	'`�0)ٷ���h�b�7	׈n�#5W_tU�Z�?�L����Z�f-��%r�b<�U8?���l%F�CY%�!�W��"�xI�D���]�-Da!)��уf=�|�<�[j�GE5�B���áJ�33�[/����I�Ւ�����i�{ �T�W��PO����azhEծ��jrk�G�
�i�	6�f�2	o���41jJ��o��f���^$�{ .2 ���n	�:��B�cA�U�}F������p[��-����ݨLU��������?2�G����0�$q�^�r��V@=�m�̑9�&HP�+F_��[�ڴ��&��>(�/P�2�>^4v�?n7WөQʂq�,,H��V��HV���pn����_ћ�k��i1�K��i�����e�����1����x[M���)vUvʔWk�H�x }21g4 �{�+&��,C7vh5�A��"��N�����f�BI"�̻v�/l$�	an�Xmm�`n�4z����q�P����ɭ��-x(M��n������m?)�ȋ<���-����
�>�IV�y��(��m IpbA��9}��F{�=x>:Z}o�+v���4t&�ŀ���9�a��RF���X�^]�f�� ��0E���<yda@Ab.gM���043�Ȗ�?
��_�rD���5Ӳ��i�����v�!	wB��^�>0 =���;hhF����FZ'`�p��ɑ�>�sm�@}g�Y�rz��:k�3� )S��`�'��6��iA.)n�uv��u�)!�#}�@H�+N��q���%G�G��o!(>�0����#�2�"��m�[/<��`�'�l��Ɔ�G깕$H��?���#|Hl��90?�l�������V�O�K���q.J���/��V��2�CQo]iwC�2��T��,VQ�t��*�a�1}Ѻ%��P���wN&$B*�6]��h3��I������L��Q{g;B�d��9�B�0�Em�-~{����8��8zn�^?�v��AMT\)����⌄�nUC�3�]�� �����eR�����}�h|�y���r�<��`�R-/�^��P�23������!)�/��YS;O���S��@Qp���v ���{,��s�ojC��S7��I�,s:�iCU�Wx!�5W�	�-�],���2vM��:ǩ�t�6���B����ЖE�������:��P0�7MR4q�����Ō)Z�=
L���E0�C"�v������|�=K����;��8����Q���f6OF��o����D4�;I��h"l�KP�
}O�MoG���v���t���0}d"'�O�?T���R'81G��=����@���a���ǶY��r}@�r�U�1�ĕ0��r�>�S*>)����Ѷ;�x����Qo��z��A���I�������+gU����{|h_S�����2���r*A#B-����:�S��� "C��aĄ@:c�z��*H��f�� H�pТ`g"4D�Ɠ�b��y�!�ˮ���ͅah��m��WRY
��1�"�wt�q����_����a(�Kϑ�-
�H~��f7C<�
� ��l�G�d��(��@L2(;���+�5H; -ôǆ���Bx /�|?F~�����l�X2ۑ���A׊��{������ٜ|�I-gi���Xɴ�3G,|�`9E�A�$}����O����d�!��3M_�KFs�zkTy@3�%\	og3����;�VĢzR���#Ё%
�������$�x�0$<n�C���b�_`�!,z�x���j��P
k/�Ɏ�?eX,J%�=���-�||�\��^-[���o<ߞ;5�a��D_J�+p!Ѐ�t�N��nC�X������R���]���5ω	z64�U��-}��ڊ��Y<�h���.��#P:!�� ���;�_T�/��9S<����_�m\MP��!�{�^�̙w�I�`\�@$2|�gBh^�zz�/�Y�\uD<��G=ʉח�������V�e���B��.
�ï�+��i��l�S���T�ӿ��&ǵ[��5)UG勌��uv�E�C�N�`RW�M|�&J���х'˟Pf,/��זq��f0&��o��l������f!>�ɘ�
4!�^��:�CQV��S�׫�Z��͋������Q�B�!@ŋ�o CG���f�5[� �~X,�3\%D ��N�4�j8��>�$Za:�F�ko�#���rޘ~�X��a�B��]�{����L*b��Pv�'l�z�bX6&"�%���>��+3Ү�2Q�\�|w-�#Tp��z~��o����L�_Vf�(��jcH����=t��)]�$�S=����Y�\��RN����cZ9n�эĠ�)��8��gg���]����ٽ�G����M�h@:�C��[�g��H��M��}�6�}�l�^��i�c�v�\}�B����t��<:����Q��x�^x�h��)l���q�k�La{�L WX�w�����e�jKyD�?�9�ځif}B����y6�lQ#v���/�}Q��gRհ4���W
�uƇں �� d>��հj�ҹ%��C�n?��