XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9�݄1l���5�U��Kĩ܅'J�,�x���+��'K�8�Eh��.�=*�a�^���:�Kw��I^��P+��������C/�yƘ��L�����{cd?�"�t��b���JEn8�?4�o�O�w�|��VL�F� q��m���ߤ���B�5�(�a����@��6��Q,�%���U��:SO2I~˙짽Z��!~�t���)*����%c#lУ	J94ok���X(ܷ�HH��6�P��k\�(�ˤ@:��N�kƕ�����11F��E��r~K����W�E�9��P����'R����f�C�>FH�A�L�Wt-���.M�U��޻<	MV�W�Z;U
91�D����,��l�&���F7��qC�4�������GQ/�h������F�ΩuB���k.YO���_A���v���!|O������'3�:����6�x�Dד������kj춨%f+G�3_Ƣ=�T�� �.���Ǝ��u8VW~?'��B���]�K��gp�c74����0��ԷW[Ў�^�$�'p����4#�^6�YDc'��;e�M�-�������4�zW�0`���H��+c�w�S��P�����I |�4�����Se���!�a��u������[�[���ub m&�
[!>MG�w�����EH+k��'԰/���U�H��V'?q�%L r-��QCl��ːˇ4xJn��B^���.�9�8�KJ�f�4��]r�S��ϊ�>Q�XlxVHYEB    b3c6    25b0�'#�eѺ�13�] ��|�aѢ'�dE�x?���-%z�.ʚ/`�뙣� ��j��9e�&��,��A�]��ktXО.�ԉ6~��Z؈���T���[��"�HL�H�z�xf�G��B"�e�m�J>�;;�c�մ���)��c�Uf��s��6���e)d�w0ۿ���n����9�t�/��f���`�iqbO\oI���|��RS��x��?$ӊ�d�m����L��M`��P3;t��H*�Dq}WtZx����������pP�����c�V�$��Ī�ǵ��?ݸ	N��~�A��<���>o4Y.�Q!'��.H�R����0�UioB�ER��:-7F���J:�9/( �����g��[<���A]���7!p���9�)Y�����G�ߺ9�u�5k�_�Ͳ�w�$X��k��"���T��E/�Ru�c�L櫎Z���(x�
7oҥs+S1d��	�TuA\��K�*2�X����aǬkm�����hD%.˛辡��vM���n� ��Ki�Y3���̮�(
��(��н�"�g��ȍ��c�x+)�/s��p�|63c�i&�1���nڂ���U&{ 1�	��N�O�MF|�n��9�;q�"W��fC����J5!��Y�Q���[��%�1������Y��� ����8m6����d�#Z*0�R�$��ⶨ*+�Hzáp�;A�s��u�^1K5K����p�>;�����ve�u�4܇�;�y85?��,h���t�Q@s:_:���nTn�S�wFa����e��`���w	��@i��:+O
���t*/��$������8]�[E2��L^�Nh;|Y�8W����һ��ɍ٤��򉪗uƂ�l0]3�t�Y��"� wY�8�Ϩ�\����Aۙ��ج�y�uᨯ��o��\O0����78�zfNeK(��/��r��
������n�6}G>q�3^��v��� ���H�`	�	��u���/�%�lKɷ�l�Y+�̀�����	�\0��7��?!4hZqq]�����"��&�9;�0��R�G�6�<5�&%��r�*�y�{��v Z;�N�&"�x\�;iHD���4ǔ��$r���N��8"�݆��Y���Ш���L2`�ޜ���H�R������u��%��I��	��C��O��TZ�[KF�y�C��2_��u�<lȯ+R��*���NM�x������������A���o��2��
1��8��j`b��������u(�.�������GjC���gB��F%?���D�aS{��{b�{�w�ԏ����&�������~n|��%�צBC\_���5�f��h�+��e��U���H����$X���ٱ�����T�#� ��ѷD4���uX�r4���񒭿�~v��gtn�Y����XRO{SۢlE�;�R�P��p���A���� �|�tT���.�`C5�V�)��.wp��X�#D�Źw:Y:�	 �r���ܭz)��%xj��F��~�Ґ {Ҩ�P怣��w�y&���a�>	�W8؉�m&j�A��̟M"
�ɼ����Oſ��=7l ��n�bI-�H�*p\��}ә"WA;Z�P���Y�>mV�L�] �*�}ex��أ�ڈ(�.�rn�`+ΕU�5oޖ�b��ti��y�=Gq�8K�A>��O��eR`�c�SC>R
����80���s�
�]����S� h���:u1L��'�ͳ�t�D�牑T���av�QɎDk���$[D�A��%��ϕ���=Q��<�N'zX�ʧq/W��"��䧃�D-/�y
�U�����>�t��`u���=zT�
��(E���Je�u�
�s�����f���"A��+͚}��X+���[�~"�f���qT�OQ�Gc��'��a�<��N�����v��Wt���l��,�EA�N���L�,> Y��=J�ս����QXn��%
���q�N'�I �q@�!z��Q�`��}M10Hɼ%�h��1݂�rAU��˶Û���^��&5oPx��pن�]�YP��y��-�-�����]ݰR�\�39�[���$G����m4�C�qS���6m��O�u����%�'��a�a�!	=[v�z��+�w�>��T�IL��R���!���˪���_-ғ	Ͱ��4�o����^���hV��x�Rɠ�v@��m�[���mc�}������4��Y���Z����b­�Z����+RE=��;1:^z�s2�妽u�A��1�L��i��F���}����
K�<�%��Կ��d`�����@�ׂ��
�8��׸|$-��0HjqV�m�F�	Jv�����.�����&��3wg��e�'�R�y�	�,��v��k��W�)���j��V����������Y�&�o9%X�ό]^��B\�!����z������nHO%�H�6V�����ʺ+���@RyV
���K�b��F����p=���F�7�˹�'��T��H,��#*�$]裯Hk�`����k:��x�U>TG��P�4*W|I���QlY����C�k����*���#�nz�J���5<"q���8�u=�u��H���W@�-ˊ�ȍ��F\��r�M��߰��L�/���g�Cr�4��S8��D(x	]�����qNw��\T��jx��1C(�i�C��[��;g���Ҟ���U����t��۰�_�	$OcT�,��12*i�������9~�|���'��^[�`�V���X'��[�lPj%��2�p23�� S�GT��\d3�%�1�t��S.�u4m甮����RS��!��=ʂ���+\�������$'��^� Ch0��W�R�7�Y:��,��h�)sd#g�`�~zh�U��?3�s;�=z���[SC������i��qCR=D�㎂텊<S੹�-����ٟYQ���p@�noH̷~B�	T�= �s��X�Wy򑄝��:�J8R�`�^I���QU������ɶ��h�SS���ܥ�(�kv<,��v-�;X���C�S ?0�ƫa���q��*�S�e2�/	��Ęa��q~m��2ݱ2|=�H�s������K�u^�{	���C��Z��V���(�/Ɲ��+4��������_�\q�I��w<��;�N�СG�t}!��#ĺ12*{u
h�Sj�<Uw�&�k�#�u��M*SM���[8G��.���ϰ� RӮLSF$ή�5�S�1DN�l.�f�>j�n�6��#�!�y=Ǩ�d2�&��E;��r�WwXC�ߑ/%&I�N3"т��7U�����0Xnk���X�h7���	}��I9&	��d�����K�!GT��p�� �yY���H�~Z��Ϝ��p����(��n�o�q�I��<���������~V��g?}�[���Uݬ�K兹��㤈A�̼�|�22�4	5l�j�j���6�'��Y��B�,N:�����~��(�!���	�6M	���dn�г����ɑ�z�&��{�����^�Np��`�$�eH�c�FI~�����NC�;�*�=$� ��=ԆjG��{����?V�ws�e�6~���.������8���5����3f2���8�F���]��z?r�g�{Cb�"��e�(��:F�h�2�EVz��������&X��R�{{G���]�&D�l��AA�a�5�zY�:{pnl�g���C۩u��-:4F�t�����6BCB�pw�#���x:X��ȥ�k��2�e@���]yj�8��+��Da��1DN,�����=*H�>�P�7Lh����=.�|�����h�͙Ǭ���0'[:.����T��)hD	�uT�h^�3��w(f�w�K��# |G�&���^���gе��V�\ֵϑ��Y?b�f3�đ>��t 5G��O��`�ݘZ������wM25*���]�,�`��>Z��[��㺝ͱFJD_��<���A}i6A�>>x�&_b��l�����p��a2��<�b�İ�u ��3�>�7����cko1VR�g3�������%fe�52�ԅg�;�ȷ�������1	�y�Z����?7�,{q����?�(G���l���PT�-�ҢF�<��X������MН����W�*������'y;̼������OtrJ8�7�������=A^�����H�C����`�q�.��qH6��Æ��g��a��-=��?��ܘZrq����bwzb�9?��>��E;�u���
x���I�WX���="�p�aPR[?tX�x&�
���j����6#6{3��;k�T(�4�L���ֲ���)��U���2���`%C�[��kX�oY��~4
Z#'��� J����.����{P(�=���!�-y�G��}�
��N��!dx� �ď4�R8���� b��]>�5r�rC�*!D=?C�nژ��T�LZ����m�6���,�X��s.+��sh�u���gva|Β�L2��C�#��!�҅�'����"A4eSq�A��=VpPg��mg0Ϧe~�]�u��̘�X�Ʊ��\�dG@�!������f�ÑԄ��;q`�LI�	fP"?j���Ñ���N��?C��z^�)���k��g���m�ݧ��H��*{C����x ���;%QQ<v��s̄��𶟢�;���� �n���
'v�zH�m/�J0
�:%�y- l��1�C;M�켍� �qM�eh��)�����y���-J6����P����n�������Ԏ�cPjn9�e��U�����`<G�+F�*�o��[Oq�(P}�����,�.TA�C�/_�/�-�.�����8%|3��6J��a����	ǌ�F�p�4=��Ō�P�RP>t�е(�/F�4�
	�����0:�h>�_��SK$�J��z�=�{�#�uu�����3�3��fX�\�f��q�8�	1?��*�fJ���p�&R�7VLA*�n�!?�SYf��f;�:\T������ޫeZֳ�s}e�螂��e� \#vC仺.Ug햐�lklW~c�����3m/U�7�[�hzx�8d�I���*��2�����i����3)s�r�7;.J�X����h�ߢ�$�0�p����ޡ���(^�k�
���8�h��ZڿbŢ��B��.�Q��VQbl�(zW��DR�-�e4��+K_���?h/�G�0�$ntCҪ����j)�(G<�ێ��E7�#8���� sx�Z�΁��O���RoI�U�0o_�Z��ę	?����X|w�!��p���KP���4�M"�M�3�����׫������'`ָ������[I2��������kA���;��1�]�ϴ���pT���,�V���X�aݧl�R����²�P�ο��%� C����/����1���zr���;���(��2�4�C�8	�I��6��9��7��,�V]��Qv)�@�i�U?�/�a{� j�{� #0��	x8O�份>���c��Y{��/�+
�Q�@b��J��9�h�/��-7E�@f���b!�MiUtD�E?Y��c�Y�|�G��m螫��hSѥu1�
�<BR��<.C�Z�C�r�I$�#\z%h�'�n�I�D�
cf`{�V�b�Yi��چ�	/6Y_m9�&����|*��*��C��h�%���a�yx2�y?A�<#� X�c[΄��֤�R��W���"��F�P���O§�18�k~�����Iك#���~ק��������Sbؐwt��{9��|�&������~egl�s��8�.����^���9�;V_h�Jk炋 vp����z�&��]k2�>���eKQ���X_���:M�΍���_v������"���J'�0��r��$l�̳N����UO�\_��y��?�t;0ϻ�4�)��ߵ�/�sl���~�N�t0���%��`w�	g83Q�Qx���?z�V��X!�{t�`���?����F��ZW��0sf6#}�[w"$� ����KjY��tq� �ږ��f4m��b9���N�T�L:l~p�����y·�]�Lq����A�vZ&Z���ҡ뇽�Ή�n<�]�S޴���;�B�G�H���Q�)>F)��!�+�(� m����=ue����C�X7^"S9x�̉����P��N�M��bT�?�"��E4��_JT��r�w�r��B�Te4��ǎN���^��0�S�'�i�QW��h���v�N;*��]n�h�c �J�
���Bq�a�eC��>z��b����F�do	�F3��d��� �״��a;@d'�#������tHW���~V�B{��1G٦
3��1�م�U�K[b���o�R��OtHq����E���݁��ض���w����9���>w�\H��z�a�Zq~��hQA���MEO���3�XD�]Z^ɎX��``%�?3j�/U�Hs_���X��Vc/���k(��R���Q_]]l��#S�ޫ0���U�^�^���<�z����uf��Β�4���=rZ�vo��)$�	?*N5�1e�L0���f�) `v�c7�(C����g5����?�Z��`SU�J�B0���B�׸(luC��I ��T���k��2F3���+�9M%�*{�'�.1�`������� �!e�%w��+�#/���I�ۏVA��b[�	��2`Ӯ���A�an.���a�G��kQC��t�y�����P�@=��״9b.�aԏ}��CN4!�7�z�6V���
~���O?4{�/�
ǗW���A��5!�Nk��</��7�	〳냾|��x8�8�v���w��
?�)�i�p�к��s_��:�\�V75��*��+���\+�d\�� ���j'�I�ťf��)U� ��v��
1�#0�.6K�$�%��8�
5�~����]��.��6
Fk��x#�H���B� ��g��G�%6���k��A���]��3���������3r��)k��)O�d�eԠ��J�?���.
ڸ�q���[rT�릔e=e���d���(ӛ�1-BMărB�4~�X�L�Aɖ9��D�pl	�Up0�*F}����^^���{�ޥ���W}�5Y^0W����d�g��M���~�'!���`��Z��o7�
Q�$�X�V��(P�$�ӫ	Yq�Y��C�Գ���*��T;��
�QJ?(h���Y�T8���G�E�.T'�o��	��9{i���������jJ�����xSiM��[�/�;LH���4�֔^3 [�ǜϬ�Hy{6��{/���h��"#w;�݆��W��w�7"b_�[�-m͓������P�v61G�eB��[f'����I���au���
���
sBp�H2�Q!��S�޲U��&9T/:�Jp���a�za8<j˓�{�I��
��tV� �Hs:�D��G��S�f!�]��������[.lXrU}C���ϣA8�؋��cwY�v p��@J#�b7T���抔V.��>#�Lit�� amF���4�k��b�h�y䘩'3gm��s�iO�C��N]�',c��R�@��s��Q�!?a/p�J�"�
5�}/�Ljg��Z���&R�T	6�|�C�V/5��2���<���nj���f lƺ]���UJ!�>̣�9�=qx!��~.�N��X,{���\��^T���Y��ʛ��ge�qC��x4I�=��!=K���@��.�٢���O�`H6O�׵�� Ag�Z�5����O�@Gid"�����`��{�Z����!�A,��s�K�^��u�k"���}O?x�����������`��$�a~�壓h�Ne ���&��������Y�$��-�k�
7ƿeKm���g��¬X����B�?�{upE��f<Q�!���g�}�o���MV�\�G�0��xk�_�uۄ^:��^�gQ�F_�)+��\�t���OW�#�L"=�P��M��W��^�y����bT	}�V��j��Z5���,E�ŏ�����D:Sq<Y�Q+jM� �;�^��II�:Ua�F��|B�$��x��h�W]0W���k�c;��fHșk4�՝���~��{�T"�� 7�wsf&�f�##� �R+��#�ԎڼI%�-Ⱦ���s��,�����׆�D����;wf:�����}�� &�̩�QV�k��}H�9�+�D6��&�+�zb����-	���5��M��}	���f��>8�[����ᕼ=��%�I�d�u�2���7�e7�~�������l� v�o0�.�!kW��&^�@M���__>Ӂi�,����c�TQ}����L8�A4�?4�mʡ�T=/p0��04��B���)���#�پ�gX晚�.k���<�P�P;s�w���V/��Y�ֆ
��D��<��{눩ܙ���"��Y���՗�[!n9���+�Є�Օ�	rf�!
���((SY���l�7>^y\��|�B�s�04�����kF��|,WXfWY�u��N�p ��
�S�v�����������,�`�<.��Eң�����Su�.�Ęd_��-�.�f��l�b���F*sYL��G�����z.�A��l9q9=+�~�^��c�1n�c����]�t�e����ʕ��W@/������=������n�E��gXe�Ȇ��0|k����+��o%�uo���s.����A�aԴ&��]�3�:Ȫ�u�q��D��_���z\*����o�y>qj �݉�?< Af���W���6�TQ���h5#e�!�_�p��F���~n���	�b�%WB�P�]�Fωz�T���B�J��Ә�H�F�x9�ߟb���"/Ɂ۵�>Hڄ�ٲw��[�r�oS
������1��p�6����oF�tHr;��Q�"Q*��b�+��O�j�~���j7 �4���Ĉ�uͷ���mL\ ݇�v���5�'����X�;i�e��6z���Ɨ���5T�L#x�|��$�ާ7!��l�c� ܻec��H��B܈���#�#��v �{p X��!E#5�t��3�#0�G�/�G%y����̲Qu��_�A{i��ꙟ�2�@XgzG�Z�wW.��b���M�V������v��y����iA�>�eUBW�'�Әb����i(ӪU����@;��$cs���T��R}�oc�>g�E��H6��a_~��7�d���a���r
aX�M�  �X�����j���ϗ�龐앧��#��F�|u�L�#���sŒQi��D��Ii�}b8o��Y\)����#�?7<z)�S�H됝L-������|gF|-���m{C
Aw�ՍZwɋ����OAXF��k��`g��u#Bx�J���~������M����G}