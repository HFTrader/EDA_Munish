XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��}�W�V�y���3���~-	�[yTHy�A�\볍w��V��U���t�֐K�FGb�.i?�::Gv,a	�{��e���Kl�+;T����w; LD��x)��5�B5��y#�}�8J�ЀwIV���D���U�����4�7ڧ�Ӗ��c�~;$y�Q`�<�xрB�:�aj�4^&Ϣ�pY:9�m�����fBx2���\�i)�m���ЬH�뮓4��T�]%�;�@������,�#4L'�#�3�w��Glλ0��*�
���wj��-fr��q*�ʼ��eG4h����*���P�Z��1�N��!�C���|D^��ƞ�����?m�X������h�;8�1٥��!y[�L���5���������|N��-��?�΋��1�V��������)���W�9�bY���nh�F7#.1��ݼ$>x���k�$fH��J|w�Yk-��YPF�4m���|�)��OI�R#G��q�8���g�d�+ڑLe"�: !2�Tb �X���q���U�SY�֗`�����f��pE��#D�{ғq�i�N���������A�W�tQ�e�<�.
N[�y�����=�I�����F���Q*j�ș3�Ǿ�Ǒ�z&"��r���L��mbM���j-0���tm�JH�D�!N�/	x2��F�?Y5oL���V��_Vڴ~?.8m��J�SF޷����/+ZU�O2����!^�B�;xDH������|l����=��Z�'�[X�K�!��4	XlxVHYEB    3b6c     e50��;8"��,�SJ��u�ó+��m��ܪEG�Ȋ�0<�Y��NFI����-[)��֦��а��p�J5�]�;�ٴ/)K���)��4Lnk�}�<it1��(�x����&9����<��Ҥ׵}jz��o�`�t&�c�H�s�����
4���B��e}��7�D�`� w����߁\w8Ť�9KT8��m�X�,(�	-��d���}�E�Ql��+#�Kq��jo�c��Ah<��'6Í`7G�HiW�na�N����jI��J�`�3�=��/ܬs2��Xy�'-oD�D%�E�;�&��i��w�J��E��џ %j?�Gg���ߗ���7&�kkf�U�"<.��������O,��ޝ9���y� ���(���q30��U(R���a��Ά��Ӟ�G���l��z�t����f����~��~�OX̭�0eY=��3�	Qs�V��]����-���:��(�4u͢AXп;�Rs.s�\���\���5�05$#��h��&o�/C���*��H���`8��x����:U��U��F�����sS��NV%����|zG�a9�B�=�NZ�O.���(�⦭{�,����zq�z�T�d�p}
�M��TC���1��m�L.Sx%���
j�=��-Rϻ܊Syc�<ʲɾ%���!�݂��aK���h������Ծ�>��r@��$���*X9E+���Y�k��� (���&�x��y��Qϴ�#���zMh�P!��^�~�`��-��ᾷW��t&=�B�.�(Aۤ	#�)��9��N��>�u�7�������Y�J�kR0�a�	���?+n�鱻�m�瑦#���}�2\|�~ �~'�R�� i�����@c�i�h���������f�FQz��0$�?B�'Y��-8�l[i� |�e]�6}?P�-�'�~�`�d���5ٰ���v\�.T���s�Sd8,\�'x!L���vw��N��(�f�A�J�6��\|@S0�=����T��;-�2y���󦊯@�U2��9"mc�U�����0�H+`��4qZ�]��nHIn���G�[�t�f���	2�F/��G��)N?gH3�-Y�!I�݇�rs���_L�z���H)ڱ%у3[�kM�+f4�C�c�xj:B��P��*�K���EĞ��z�@x��E3����Kq/ q��:?��ʀ����/�����\��Y���]g痰ye�t�.Z����TV{�rgK60����(�H��(�30Ҵ"(�W���"�cyk_��Y�?a�-�m�r)M�7b�F$�[����'��DO�� z���U�&.��Iډ��s�����#~H2��_���x)�J/�H�:>}��w=�"6��H*�|$3)�x��Ad���M��3zV���ҋ<��d��Ӄ(6M��B>��n�@n�o�V5��*�&+�9*�`FjXi�?�s�&<&M� �I�vi��5S����"{ZF-?�9�3�$g�D��uZp$&űK�í��f7�׃-c7D�p����-˒��X��~�'�:�?Y���e��L�Q�w�
�0�!�9n�|����w����i��S_���	��w\{x*D�t��R��>�scc��$��5pzM�5�>����1��H%=Y���$��&?�S���96d�(nѽ�t{)9���nJ�>'��:��=F��x�
99�=TK��or��@�Q����|���njqU�ح���~ˡ�Hϳ��Q�n�;@�����a���c���cB���]�ˁ��2���h�;W�r�&A.��$�xOɼ@����Lq_]Գ�ϪAW]E�Š���P��{��\h|����Q���/����)�I�os�#�ox|v�{L�lR���dڇD#%�nn���<�M9��=CPH)k������7Dx*]���%DRt�n���;�(�٪>-rDWU����}����ý@XY���i�%UE+j��B+��éx�U+rq0�S��)�<�f��w�P ���R����<#)SN��R[�F���n`|�0�4���D0Bm�� (c�{b Í��{�g�DD�3��Zs��E�L=�7�3T����"�@�D����p	�5{�� 2��ޑv��b��
�w���	�#ڝ����)É2?�0�U��$�8U�-p[�a�[���R��!�&�$+��&�?}�C&���R��E�d�m�����h��F�Ǧ\��^J_�٥��M�je�`Ure���ǒ�t�N*-Y.��#>�[TF��;�ۦ7�3i��b�;$?o���e�[ U0ja��)xr߻Q+��:�;ih��ޤu�J�� �J����v�!��DH[���\�a���k�Ye��|ik�r?���|?�K�΀��ńӕ1u��2����Y�4�M�Z%��7���B�И`M�8:�������j(#M��QaL��$Tr�(io����Q�M����lض�ˮ��=��11K���?�U�#�_�pc�;��Ly4�B0�BJSD�ۯ�E�A"!�1���紤�c̟�:*�s��7�<����w>�7����`�bT��t�N��˴�4��P�n�f�<SP������c�QA�L�'d�J��Rrcp�$`�����������9L�T6��3x�@4.e��1Z��C�Y+2z�K��ύ')ꇜZh��9j�����g2��?��|���-#ظ�ӣd������	Hfc��m�AT4	� �G�o�f	��-gT,
��+k�#Z���U��^R]?���/V*�z��#����� r�ڒI�Vd��3�3~�2X�K�J��8�x#��]K�<�H��2�/S������E��6ޮ�OE���2�����'�ݴ��B�̞(q1�T��V�)L�K=ˊ�.3�ޡ���S7��{r9�]�#�qM�m��Ug�XZ^�7�7n��iSl�L2��p���cpآ���W�
�
2$��j�k�'���w��y&Ϳi}L�y�胩Y^�V1����q�>�!� ��,���rG����	�/%��Q/���s��j��,,�o֪��{�ˍV���ԉ���� ��5Cت���`B��i�ۇu ����X3����A��	�>�IzϏ���2�_�CY���12I��b�G-�v��[ ��U�t���)�B�s�;�Y3 K�l�ǀ �r���mq�MD��2����a*�VS՗�>F�<��ͷ!X����} 9B�aJ����$/����MyG����@dY�n{rx���)Z�~h�ꮤ�U�V�ò#=�5 l�O�`_{��="���/�]�f�.KɃ��g�(��d���A L(_�h�Ӯ��ں	�p�W��š��y��I�rAI�=Rҹ��VsU�9P#֞�_i)�{��" ��5Z|�N��������cn����J�Z��ًE"r�-%�"�����(b�޹K&�aGh[���=>�a���cpڋ�6���3نE��	 Ɛ'�Ť�?t!���e���M!��mT��i�/�z("����1���?0	�f�Z)nޜiM�<e��$sZP�B�'�aq[I����Ϲ6[�]�m=SU�r�+�?c�'��,G��IO�d�!��
=����� 