XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����wE9P�����U��}�d|����u[+��@��N�+i�$��D[]/o�H�C\����,̫����C��uw �e��ȳ7�8�Ů"�t���u��j����g�/ᓠ�iM��`w0����OX�]��v5�`I��7�Lϔ�M�)�r�	gv���+�q]������r��k�ݦ��J8d>�]���g;~$�����5m�V����L����3N�� gx��Yɔ%x�]� ����=�m��i�P� ���&eeC1}^���ky������csd�ts�-~7M���]�%��e������PRM޾og �{�x!��݅9����i�A��%u̱߮�Ru��+�4�8�� )�)�#����1X݀"t'?�CNj⥳A+���L�Ӵ{�K�db�Hhn��]��a�碻���@=t��jhW���;�"�����z����^���Y�D�,��+1L.ao�nG�J��	��+��x�ꏫ���Kme��)�H�x��ۧe"�,��[5�g��&�C(���?�#0V/T��X��0.Fl���Ѫ�~�����!8I~R��1�o����c�����9]$���4�Mo�S�f�m��%n��<(C�����$��b�����a�M��i���N��V{���Ru��<k���@�m?���H"C�x�Kꍆ�J���DB�aifs��o.�@V�h�������w��\������4`�Ñc�����ƫ�/�ɶXlxVHYEB    2577     a70���^l��ˎ���HF@��f��j�Q3b�F��}�i��>v�E!}�H��[=�7`�4�����ٱ:2��AY�:��;�$Q�*0_U8R������I�kp�\���3����X�/p��j�K<�>������������	��+-&�=��-����"^�m��u�B)��9uo�]&�wC�)6�2[��I �@��r)FG�F쬸�>57�@��Vݣ����5`>�V؊�L� {����&��)6"d���rX��E�c^��ɄsoΜa}�'�,�F�t�.�{��凃r���S�V5�S���Uт��(�ShC���JQ��T�y��z�$Q|��{��|�M�i��X=���D#��G�@Q�(ue�i���P��^�^�.��B�m%.�J�L�e��~g	5�r��U��AP�z��⸀�
ʆ���Ub��E��(0�q��w��?{�"���.̈q` �#Ȭ�̩�y�Fq̶.�8��6��2f�R%_��Q��N����`ۍ	���hD�22g�*;B�ʖ����ݨm�V-�[�~^Bu����� �jn�x�Q����Z;i	a��\�F#�orRq�Ü�O������B���#� 6�c�H=�����X��"{�t�љ�QF.�H�^���Y�4j ē��z�D��G+Kn��F��1�^���=K�)�O+m��f�L�6	���q����xw� ���#�X�-T�+����F����M�:��1��Y�+����KZ;�,&D�T�eɨE�F��{ܔZ?[�q�8�|{QM���0�_��\K��\�\#��n�!���B)��� T��"Q�^űM�B^Գ7�rɝ�J���ĥ��Rӎo}����� G��L��U�M6Dy���\{��\=��xUx�L �LU���U(�T�`A��T=;�j�}F~��d����Lse�|&e�Ͼڪ��O��l�`�h�9�d�Rg�E��z���F�}��m�G��<VGxd�F��0��N���>G�ie��8��om6��d����M?�7E`w.G`�Ә�\�<�|O#؉	�<Z�����l���m��Cl��k"	��O�?������"� �6�ugӱ���������s� ����{�9BK�S��]�ɚ679���+O*/��/E����o���C4�[H�X?���1��Ǆ[�@�<2�E��\-$��������V��<�J�1��}�:q1�����aF�����kf�ʗp6'��P��ǻt��E,�_kiF�:�vJ�$��׶��s�O��n@?������0z���ÛU����#x	�Up��;*��y����P!���:�_gU9X�GW����#]�hD!���������	�Xv@�Ll�=P�c�`;g�L�*)$�'���['�%��;���(�2x13޹O&-��G�=ꖀ��_������m�*I9���_�;�f%`����_�	�v��W�z;�R�I�ξӭq�L#lgaB��@��k�q�@`S���M�����H�n!���\�uP6�S(��$�v�5�2�
�0����46��tē�ѧ��:$����#u}#���"�s8�����R���$�w�gHY�U%��|��0 �Ap�rg�D�$Iٷԟ��H�c��W?��V�e�Vj�O7ԲyM��� �?��0��|��˓a�G��K7��p�{��O�SH���Ȩ|�!����-�����=^������T3�?g�+�W(c����TR^�I�ǚ�\\��B=<�%{��h�.{V}�x	��qی�Ͷ���)s%���i��ڂ߯q����A	_��do*�	�u�#p�� 1���~3Z-�Zr/+-Rʩ��uo���iƩ�a��#a�/lg�V20Y80�Z���pUd�p�{�eS3�O� ��mi�Ȓas,��O���,��Y�vb7}�R?�	�-��$�Y���a�±y<rX�_,�K���h~g̍ E�O��e��������l5�T�V�|�rE�)�`�6�g���nx���� �
�T�1�7�^�M�Ԛ�l�Hbk�����Ɪ���g����r�UoK�3�c;P���שNLG3���	�7b:����4���V���ݻ��|��p�����B�ԛ���B���a���&�����,�����RPI��~��}��qj�i�ְ~�~��F�A�h����d���)��T-E��7y!�#�Mt?61x�� �O�T�R���ؼ���m�ԗ��͌g�J��i�u:�����Ip|�b��L�Ǿ���%5��:�
����Pη���p4	翙�����8xa��B*0C3�;Y���	ծ4�pa��5J��]կ�"��g��I��!u ��!H*��}&7�<|�%O,0�
��wL%��n��T4�P{:r���Rӝ(�T�4�@� �\`�} �i�r�}�
����Ǵ�!����K���#|�9Uz�"����V�啯(E��ɘ�[������*�/����5�'7�QL&�l j	�F���d���'k�m���p~�>Ť�P�q2Nc/�6'�����5 >�{$ۭfB�I�{i�7���������s����p�X����@