XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����x�+�=���[��6�������틭���C3��O��S�a�yBa�U*�������a?R�Vj~�H˯���_�FůcįJ�����1��F�X�q�����Y��Y��Z� ��|�!Y�>��bo��d�+��a��7�Z�5��:c:h��S�ì����M�bK2��88~)��6<r����OW�� �,�VY�H���W�$�÷�r���h�@������ߪF��%%*���o�J�m�����lnv)��>��AG+��q+R�C��h��_<�j�J�Ŭ7� 68�u���O�Z�W�L}�� �3#J�_�p�h1����l��-�q� S�����`�$��&h�aG|����!@Tuh:�2x���{`��������dx�Rǘ��k�Ul��_���Y��3n3�kn�HG	�®�'�����`:h(Z�dd�����qd-.#~�1<��?����� ��6��(�1����x �f�,0��8)�$���M�n]+AD��T}>�f^�j������eZ��|%AfJ���Eez��B���t}z�ʩ5�`�׷1e�@�[����g!��=����y��̬�8���䕵 v¨ �b������,�O(g梸��ы^��T� ���m�����7=�� A�tfMd��-��P$#��"b*�@e�7i IY�������Ȱ:O�ر��2P6Ñ�s�;R�P��Sރ�;J.��4Ըn����Oܞ�a��	�m�XlxVHYEB    b8a6    1ac0�N�4�=8��l[��S#�X�`e��4��P��;xKeR�z.�"�<ћ���3�^aXa%�V	���y��l!�,��Q:?WpB�ñP?-#r7M���R���>2�<�c]d=܉��+Om���Er�8�(��퇈Či\���+���%������P�^���*��w7GUڔ�Qw:��C1�CJ�Q��~�2���h�#+u�������T�s��2NX3H���&�O\9�a#so̹�#J��Z��k*�Y}H�0��g��B�B�۩�Ԥ�wzi(�f�-8͠�O���������h�B�|5�N��;)A�r7-���$�N�ї���q�N�3�Fh���4�M�������Զ'd��������ѵ����
������mbEl�?Dee�Qe],�i|Ӎ��P����Y���VI�f!��I�;��0M��D��
U��.����Cw=�+����h���ft�Y�n[�$�Q{}=S�����z���*|\P+����vss��D�f��+נ�nYgQ.JB9�j�n�:��x׭D��o��� ӊ!X�87�vdm��hF��(05?!�L����������%��Vf��^?���/{@LwG�\�܁�X �+W %ϋ�Ĉ|~�$g	^���mOk�>%@r�e�1z��Y,)�yKϥ39�^�-My�f)��0{:*��ܮ��}_���~���[�J �Y���Jk���]p̪zå��ԏ���Q9�]/~�'j�z�����QKX�l�-�^γ���獐6�����YliTZ�:�Zo��?��<@)M�d���L<|L�0HF��G`o��⌄P����ͶpQPa�f\Kb?.׀ � FL�Q���>���:��%1��Y���X9_T��,����i>��(̍�b���'E���T^�b"d,T/�]�,�`��3rz�c�:�3`�le��U?O��<�&ϦchS6�p�%�y�m�"3���+��Cą	���Ľ���t��Y����̚4����0����џ�y�!6&H���;�s�By�M`j.�gf�P�D1�S� �_+9^�)zl��S<]30���r���f�:{�3h�� ��e�Һ$��ߞY�T/����)y�3v�%�0����V�\�g���=S[e'���0��u��O`������`�ڷIWP��d���]}�.w��##+z�Ұ�[3��"���D��\�i��� V0�t�"b�"�����q����9-Bj������Z���k�� ���:U"��*f�$�g����(�Oɏ�ך?�������c�S��v�!�/bS�*\^|=hLbZ"����esY`��Dh��.��#Bo��͒�;W�*w�r�����H0]�f�H
��b]q!��@-9�2�H�,{�2�,�Ą��i���:h;ݴ��A�OX�x�H2j36�4|���B���0�����e$��š7��tw`�+]DrF���<��<t����C�[�hVF�Z�dR ����"M&�w�*�I	TU_ΩK�	����V�R��'�L���c��s��;�o����)'J����0%[~w W9%�3�h5-���t#���W49=޸�x����R���R�F��\2g1<�qA�V���NKA5��׋Wӎ~˧��SJvW�J�Y�X:a�.}��6o��S�B7C�h�h�K~Ne���Vx����ʼ^�q{g�?@�4�&�d�y�wZI��y7���R-(�֋��#��H���t���)E��as��c������+��N�7�k���V�y�������s�������,��O�1��� <�<�rYg�	ߐflh�:���_ǲ�M ����_��7r�b�PkZ�yV��Č`��NJXIb�a]�Y��ɜ	�������W��}��?zXP�M����p��T��8M��S9�0�	(���-�q��r�!�R�ǄZ�S�6]���F�-��<�LYF��j��UV�6u|v޺
����4#���P�����kϳ�E�������r{={८�r�T����׉����b�]����ds�������'{�Kb˫Rѡ�j�!���B�.։k��뗌�%���ܱX.Zʮ��l� 2�a��V��A���M�dǳ��ʍ�V�_m}e��d�@�1@�_�� �.��ғ�?v��H���_Zd���y�^~�0���g9����z��+9+(�h�� �d`�����=�nG��E8C�k܃	'�:����W$:δ�Y��ߩ��?d"�����?��E�\�т�J�/8A(�m��H�:�����W�ʒV�Z�r,D!��׵��*Ƴ��"�F ��u�mVٱ��Fu�į	���3|��vn����u0�|J���P>Ʋ���ы����n]#� Hg2 }8"��MVG�3�~k��N<�xǎul�i̋N� �~D��Sߎ����N
e-�� �~�i �sw։;!v�.LsAhiq�K�R���GnG�+͇K]�G���t��}�:�1:*��H���\��W9"�7��A�!*�"�������g��G�{�0cp$ʴ>���"��RE`�,�@^'���*�s�k�ZIȔ'a��
Y�v_���"�-����@
�a#�	L�X	�)��^a��7&I.c�sSOd�x����~�!|�xi�������0�{͉�5����4C������#����(�>�l��#Tx�]a��j
�����\ZR��Ք��ޣ�F����˂�N�^O϶Ǚ}�����m����+Y�b�D&cBI����؃d���t�`7���ֳKƢ��I]�-�h�j'��MC��&�$̃`$�w�r�{�ںK�?��F����OA��.�8Č?g8�l��)���B�+�;r���N�F�xe�v��Z�%���0Z���A�M:H�~y��|�Q ?6�V�t�oR�ؐ_�s�d?��d���yfNe|��5��)�qL�}(���yw���;�ؽ��RNEq��DQ�

�J���t⍍ix{�Yq�|	>A�ԝ� �)Zj��?���Q��؜i�ڳ�T����Q �xF?��ҳĤ���]�d�%J����f;�*M�W��Վ<��B)a	O������+��u����=zgw~^�np�s����������'g��'1W��<i<� `� #��6HS��ɖQ�z�Ӏ�P.c�_��ɋ�oV���Y�|�e���jD�꣹)(�kF	f�dӱS*Pί�?WةҨe��&[$��i��N�l#ЕB��Q�]�Gn9��Hm�?��C�����l�؇�鶊�.9��nT6/�U�W*�<�a� �}��ˎ�Q�]]5�jk8I�j::��������m�����$R�)�
vLt��i.+�R�ow�W�q���T������$�V�!q�>��L3.8Q^/$���]�	�֡�[�ڠk?�Zg�3���/7&��&Rj���_��6�ӑ?~��Z
���qA��)+8�ˏ����5j��-�/Lyc�Dgq��;L��lmS�,��
�ؿ�������x���k^��^_NN+DM��l�"��xNg�3�𾚦��VÞf&"fx���ۦ���D�R?�� 2h�����>�x�.M8�R~��,�|z���$��D ��eR!3rc������
���'� �c���a V�ﮟ�\LqY���@�[ڹ6��y�A�9b����\Z]�V0�V�xd�8 �X�.��Zn����/�T���à��Y7�$���)
�淹S*��U�k ��+S(4�q.&6pp�P��q�?��
׀>�M�j����C��1�Q��ty��qʿ�w)�rE�)) t��U}�z��1����3fJ!.L�5ڏt-3"�\ղ�1�� 
��z�ֈ���{TH*����K�4��ME�i�ɇR_�ӄ�g1��<��J�,�/ם�y�F?Ϡ�0(����Of�"�����!)�E��;���)[�����@�Zb�6�h�^��k|	~��K��h����i|��Z�$YM��qˣpSwSg�O#��w���*��h[�vL�xXR����ň(���u�����[\b�z�=�"�O=�,� ����<�7-�,��u�8h�c7�a�Ɩ+�ds8�����~@��N�S�>ս�>��s�Ee�b�H����INI�E"B��-�1�b��\�<������d��V��բ`�}ђz��8��B
�u�������헼�����ȉ_n�!�MQ2@<�˜��<o��Jur9���
`�ګ	@Z ���삭�̞)�?<I�di}��H{q���2	�Փ�p�u�Q�N�'eN��ѤI�F�M�F�q;]����b5��D��;�V�7�,|H���Aj�"��O<#����9�*��\J�H1�KFZ ǰW"'):��{.����[�4��L�9? ` �Ψ=�wd�FV��p+���y�I���{E6�3I|�K� .H��'#v�����Դ�F�k�+Ƈ�5��74^��;#W��D8����X#_�\*��fⴑ�}��P�CR؝����� ������o՜����%1��%�����UY��
�&�gv�^���I�U��[�]Ns;��m�N�+��/�xU���;x/���CW	6�a��$��T@���: NE���`�M�څ�_"f�T���8x�����I��p���P��Q.�����B�߈���g��-h�a#�!E.ʊ� @`����q�λ�Pd�`ډU�K��_�J;���A]5Y�p�,���3~(�\E��A\���1�O��
�Ε>$4�t��;A�����ȩ�����UI�:��s����or;d�g�2J5�-X�����_4	B�s�),w��
���b��2�\3���!�N+�Y���6��Ϙ� ���dl@���1V�������2��GU:�p����#�!_�Xxjf�omx�?w�-�����щ�xK+��9�nIв�g�nٕ�Nr�ZY��Cr�S���iy�Z�p%�A6k�@h��n��F�;���wY�]�h�U"� 2x��}Ԟ�*2|:њ�p��H!"M�9/L���~�ͅ�IP���*n��*~S���r5 =��z켚4�"���������ט,�\I��]V3�fZ:^� ߝߝ7�1<��!]��@��U���A'��E�Bu�M�fX�Sm���������aّ��e3�ͷ9_3����P�Cδ���	�i.@����7[�HK���?�?E6e����G$�Tԏ�
=���J���������sl��q���{�K`�)4-i�3maSeM�gx"'2�b��)�=��2C�L��ۂ�!�dhb��lh�6�˟:�"��������?Ȓ��~��U]W.�\fqF�?�.������&�6�X `ыCn��7&��o,��H��()��W�]����g�,4�k�K��������z�o��Z� ��(_��*�C:�V���=u���h+�M�"}!@GI' b���8Rs@�(����{�����w��!����Z����b꠼+1�ˣ6��&	�3{���/f8̖w����#B�N�}��q�Lv?���&������R=��s��`����>����v����#���}�����H&S.Ը[s�-[��#�Á��Z'��*z�����g�JBI�_5���$㓪!w��$������ ���ɠԶG��v�����LN �"�\tw��=b��wk�vL*v��qN�O�V#���I~�Ȼm��]R�%�d��X߹��?�Flh�Dm`�-�F,��:���h�m�>�"u����E��
v�R�yEac�7�fy7�?��3k,*�k��Ͱw�]���������"Ⱥ�Ikl������)C��������<F�|���=-޳�V��2��y�*7�TԔ���|�H�8)�9�^F`)ܶ��L����|��2O��]��q���������z�����a��)�R�x	WR����Ɏr�����)�z��x~���-�et�0���FA�B���Ӱ��һv>�����e��P"�N�&���X���U\��7���s~.Zg���L�?ߞc	���}���,{P^�,p��Y��/WJ쥆T�u���v]�.���|d���[0Iﳑ%�P����>+Z�\J.P޸*�d@23�<��s �x"d\n���4��Wx����!p���L'��>�:-��U$CF������b�s)��'HQq�G\��^#n|�E�]��O=�vm1WH�'u�9��"\��p���b��R�pQ%��$��)}Pxj%0�\��G�$ή��(�B�!{�3]H�|D|�;/:���&�KoPx�$Y\�I:^�L0��ZQ�Y3vT�p)�e�lcА�#�`w�Gז��C�&���c����!;��1GNV��t�b��A����4�Tl:������guv��%ƫ�-W��?��"��F�Y���{Qc� �yT��a,��EF�������4�߾�r�o�(��u�"��g����Qz��E��b��2TL��:z��-����e+�¤������ѡ����L��[:�jqW2>�~���j�5�Yw?��̦��Z�ό�^	��&Ɋ�aE/D�E�~O&���#@i,�y|���3��ݐ ��+r�n���*��^�u�V��8e���7����������a�t	�����Yu����^R�Y;RY&69������ɵ�泻^�n��q����]��j:+�r�^���2L����LÎT�