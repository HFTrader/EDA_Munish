XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\�G��_���'/`>�E���<&~P<$����9�дM��! �P��+�8`p�������$ ����_k���a,(�s""n��#���5~�E�	�gQ��qZ�����В�:V�Qm�̎M��`�e/9�&��#{jL+�)�Q4E7�|��ؤU�?�]CY1x��i�	+3 �.�V ������J���`7]
]��W{�X/9�j&����62��Tk���[���x�.�$��/v���ʤ:O�&W��'	� j�73V�!�1J*\���	��S"W	�?A$��XI\�_o��oM�ѷ��ݟ�*U��� #zx|7�1�儢��3�S`�<�{�;)�:��	e�/f}m����l��Gёd��(���7��rY
��jg���M95F�;�BG�c���S$Ow��o�� �+O�s��׆k��Z
������?j/����7�'�|�|f��!�Z��}�c�UDu����Ho�<��A���m��_�{l@��^�D� ]�����4���8\q�|��0�����Nu�KB���qh����ۢ b+���٠�L��ѐx5��U.?t�H��ȡ�bw9�4���mњ�	'D�Du|�:EO�cVK��Y��lcD��
��r�h@�%re��w�n��v�wJ��N2���'�8���2Z�|��X���Jvϡ4��/?S��"1\v$J.O� P�Ҙ��y����T�r���s�`БӢo�������DH�D�B�s~O9�UQ�U�PexXlxVHYEB    3099     c405q\��(|�xg����gJ��6g)H='gۚ�B? tJ��/?� �s&�ҥ@`��^�M}�7"e���D�`OR:$ە�x�_�e,{�՞��4�C-�X���v�H�VE�m(�g����`��(�O��]Y�����&C�Z�O ᇇ��H(�P���-Bj sJ���c�ɭq��L\��n|�{�Z���\§r���},R9h�Lo�y��(M�+H�Xa�w�7�ೢoX�7��
�A�$�A����[�����~Ijz3-��ק�^�,��oyb�?t���
���W�_w�62���8��#FsB]
t� UKd!�$�mRm��F�I���ĤJ���e�g~+"m�]Z��ԏZ�^���4����Î2$0���l�����C��J#��e�Le��n<X�2G�����pЋ�0���%�����RN%��c����53��/>�.�G���`��,�Pc��v��lH�����E3��'E�` {���E�/����Sya�F�dٰ��"�p(#]�z��)�i�qr(�QN��M�H}�@� �J�����*|���g>	)W�����1�J�����O������u���5q��\��FLc���|��m�hJ�������I?�䑰��iK�W�2;��a^ZtS@g;��oaOW�ԜHp��x�Nf�*�q�,��w��F �Δ��_�r��"�V;�?�X�������.?H�E�莬<�G��lВ"����RD�f'u4w(dQ�9� ]<8Ƽ���e=�@�h��;��V�`dCRQ5�"C��LЍ��<���/�)},s��9��@�n��?�^��GH7�?'�-���r��IY�'��Y��u4�㎍d8,�y�X'�Q-H�I����
"Y����)� �%+^�8�Q������Q�����-��46��1?S	E��Bt��Q(�Kq�C���I���oɫ(�L_C����=��Ð<��7����	$HDE���y�|�;I�� x� �D��ƍ�@�7*R����qT�r�lv̻�(���"���k�z�44�Q���4�{�_����Jɋ�L��.�7�m ���f��2�א�ݢ�g5I(e��Vc����;$e�ڴ	R_m@��Ǥ�GX8�+��S�I8]Z��F0)%?R-�Zڳ;�<�w1إ��(�lyM��ڏ�{�1w��w�嗽!������B�C�Y|fe��>NJ����3x�J�r]��M�LA�l�ץ��I���ѵ,W?��z�Br�e�_�nQ�[�pA�$0x����	[��͋����yYu�;�)zI�Q�E�5�_�N���[�&��U�N0C�\�Q�����tb-�C���@����G1ݎ9�6"�7)][���`Zrmtჹ�U(Q��� ^i(��*,.)f�r�~������I�-�00�ē�����k�wȈ��F��.�!ڶ�_1����d�
��U�Y�7Ľ��A~���c���;��c9��j3,���;�iJDI(�U��ߚ��|������ub�F�S�� �#iz*dp�aP!rN�#��H�MT{#��7� �{����f�7�t �jHl�Hŧ���&���V�6�D�f�����vq�AIώ)/u�c���)���*l�6������g\��0e�4+[�g�/r���'c���{���ˣ�4�'9r UB���Ɓ����ڬS�)?��~�����ibFPH�w�X���֜IhͲ<r��|u@�J'�k����	4r���~�k�aG�{�*��R��:�Xs76L;
.�?�����0�~S��%����]�J5�F�[��_{��Q@�zBi*���E��߸�\�*���w揫��+H/h�I�Rɦ=L��6� �������܆�R�J˜E���E:	i�o��!��ֺ��r��o�h���L�8f1���,���y�C�����LS#5�?��m_U�ϾW6;�lH|�\'���kC�j:��݄j�԰��,����DN������ke��N�2ɴ84��_�8�۝�^�.���,��ץ7\�����\hn����&� ���u�.ة��^S�xT���[d�È���j9Og����oկ(���Ct�E���]ZO��-��.�T �ex�Q�73����|8��MC�̣m��rqMz��ҕȦ�8Y���͐��S#��A�q��J	K�8�AR)��7W$w�-�>���d�1�#v��y��l�-D�^f���A�� ��f?�Ji'a� A��5��[1��0N��n���~���WRK�d�!{pj7m1�g7�c"�:a5���h��.T���:�����3���x*o�QH��a-�˾(�2�\O`S���
v��m!i���e���k�
;(���z�
�� �\�nW�
�ja���(�:�9�+&�B�Ի�v�;���=���p|��#��8��qLXx!{i�J���'��Oy��U�-�6�Zt%��iF�E��x]><:�;i���O|��[�{���c) �Q��M���`�eu��`h�Ő��f.���m6v��-�̜�@K�K�+Ƿ/�#2-r&�v�a�
�6������[�gk<�T@�-=��HH�493a
Q|���ێ|XN�������J�Ilz(���Yq�и���K�C��\6@�9��Y*�Ӡ{A{$�5y��@3�����!�+��������w���Cc�V���V�ߘ��#�2���*-tG�>�p��B*��������B�b�k�u4CLT�G��8��������(��>���?�{���㺢"�c�����%)��ᮈq$,���Ϭ���a�ɣ]�.$��z��Br�>�����K�
i%�_'���F������rR{�k� ���R>ڤ G�
p��u\[�	c\�э.D��&Jx���zm5�JJ����0�r
c0�Ѝ2��_(*����!e�J1ϝ_�Wh�4�J��=��L�&c*\$e���ɆR���cňl��f���e^0��\wjQEoi�Q�\�όn�y� �����Uqۻ�t(�Yv<�����}�d�)�2�Er)��2(jK�4�b�z+K'�H��D�F^~��M