XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����G~0�B"!�9��~s�Y1V0r%EV�)�����_��S�T��֓���&/��֍W��O��u�x�I��-����OeU� �|<q���E����q��C���O��04ke��2eL��C�n�{���i��km⍟�
�P��܈q!�����3f��x��.GA��U�0.��L��O��n����B�?mkj�V2 `5�~�d�>�+�tPE�?�N�-
6:�(a�.=�IW���s��R���Y ���ÈҴqwJ�BY���Li����qL�H�4ܜ�n�-������L���}�K	����Wa,���6O7� �؍���/8�l�!D�����
�A�������?����?�4��Ѽ/�߭Ӏwy*j����n�s'֖�y��4Z-��MY; (��{��<Z��F������t+>o��<��)��ZY��Xn�h�o�-c�?�Z�k���@���5$J���2�u�s�X��ikt�}�p����BN8F�7��#|� h��3a����������Z�΄py�_:ݚd��������o{�
���Hb�&�_���}��{_�u�,�*4�?dΥSG���ȊS�� �"��'�2'�М��0�f7O?;���`e1�6���G���؈l  �j�K����W���{T����FX��-`DuJB��2Q��ND���<��h��/�����z(A������qԢB�^�;�f�*��۩&��XlxVHYEB    549f    1060
�i���@o���U�<]�͈��1ZGVW�����ͣ��N�����"� '�E��O�������~� !��j�}��z4��J��5	�e[z�zo��J[�+E�"�u����/9�WM*q�6�@�x��z�̐�AnS�V^��nR����8=#C�C������Q&V�s�Ȏ
�8ʻ���ޥ3i{�}���u� ѩG����B���Ju�����Tn��t�'>�i��8&pw������-	̇��N�,�<�H������o/NƔ��ā\���$ ��ϐ\a�� �h"�0�0;��8�0 :l������Z���I�΅'�T^SՉ+����Jp��,2fXv�L���%�t�Ld�sp����[(�CG�?��W�Tu�AA�%�5�5�m��ܷ<�j7Ԇ6s�0N�r��6:�@�|��T�}'<�*��b��p�I��[���'���Q�N{aNi�q(0�-�i���6���!�$�T�����2�"&O=q��� ��!��Q��6MHz�z�G�����4�����J'Ef,K�|�DT�� ���o`V�PPt\��)U<�%��x�)cQ �euL�Q�ڷj����5��� �Xì�`̻���%��P����!�>�K�.i�N���l�2J>�>�ؓ���v7�kw�����P�ϋ������M�fZ<(g��M�J�¡9F�PN�+]1���uq�&�gk���Y�8�	G�?�~`[>��Ã�7��
:l�8���v^��� �цõs]�@�S���eD�,s�A���OcҴ�N�S�ZZQ�_E�=��k���eM�C�� ���)y�'���w��0���S�(W$�F5@�Ko�� h0xJfK7���;��%����C3�DC<�U��7�趉��W&Ij1���bP+1Q�y< �/�.15�[��HW4�$cO�:$v�XS���`x!%Y�cM��rЫ���à?��E]I/d��:�
��&=����ޫ�m����bF��i2�i�aс�m?�e��}���޹e�O�pfL;0a�G�+�k�<f~`76΁kr@LK�d��u�ԅ3a��Z���� �����G����R՟��'�Ɇǈ
���TZ⅞��O��9`y�"���!�O7���De�^L���gq�ά�K�5�c�U�����?�r�ɺ^e�]8�#�M��y;D���Wɵ���.kQ?�;�ﬞ�%S�-����`�B]��߀,|t�9
�>[yG�9����EH��
�x2}U�04����|���g��&��G�W���n%��ĉ��r"\W�N]9⇇����hV-E�_}��=.�!+���8����iQU�Ocs�|B�tRM1�o�����6�N���-O6��5��@�$B{�N�y�xRG̕#��o�H24�0^����N����K�jq�r�p��~
t�Ax�QH\�����N�~�D_L^���� �{^٘�8`h6�e�|�~����c�/������g���\z�����ض�`�T&BS��\��e�q%A!��XD4��Kު���:�q�I��4�ZT��o<��	'�B�+�t��@�����Z���&�=������d�Z0��؀�â���oG��7�]i������t<��E����z�#�\�Tfц�
.}�u���ޅ��������|�� �M�}�������u�!���),)�2��p�.�!�8�,4�Q����25�!;�qjS�q��8��/aΆ���Bw�W����o^]*]���ѱ�ꈃE�)u��[=]�}��8���j}���-��L
)E���� 		����ǘ��~�Ep?�[K�@W���I��8F'e{_�H<1��b��r�.k��:�C���p�ܹCRepo���*$�xkP赈������ہ �~�$wڝ�k�W)�`[Q�è`v_�`:����U~ocJ=߫��ƒ}$'}uZ�%���>�	2���L�0A��;3���'Aγ����>C���g���߇�L�������v��Jy�By�-��J������⠘s˹����e��_��-mka�1+�{�pYݓ0��F�u*f��B���/ꥥ�q��Yj"郤�ŧ�(�"��L]���|<e�N�n���}�K�b�$5:�#y��>�������U�d�*|�LH���~BH	G�C���r��	��b��Ŷ2�V�n��Y�`� �Y.'ȭ�(2��=�ނ��Q���2E���?�bÏn*����<���Yc��F�mB��_��9��Ɓ�����I���J����S������uz.A6�$�3�bP��{�ϐ7ڽ6�Β�=Q�����t�����<hP��R;��!��ze(��z�Z=����4�ŏ���>�=�H��!ٹ��8�#��2%��!pE�ĝ���OܯՒ��h����M�U��l���L�~A��֛r�I׶A�)��:Uv�0��!r/����/C�}v�B�gc�B��jm4a�#b��W�i)��p#փ�U��o��C��9�6��N�]��wV����h@%����l���X����6A����n�gG�N��xぼ� �� ��F7*�����K�6k=1�1�r���h�����I������z�3�
i��;����2~���LlUL�@�_�<� �*�w��r��`�9*{R`�%�%_�� ��%["���j����z��e�(M[m��
��7�N458EUQ<���T�V��t����4�V����&lP����2��u���V�g]?7 Ǡ	4u��z�a�Oq��%�M�.g�	��t��K<�I�v�"�C<�_Ίd�Xe�{�
��^'�D`~�� !�)��i�Jn�*B��'_n��N�Q#��-���^lb �q�HY�^�\��2��,�둝X#��>[�����W�D��"NzU�D�YS�1�S;1��WV_�X
,�ǰ�$򅡣���h�6�O�I�:��*W�_#�UƤ��������ȋ���)�4�!�y,O�(�����t?j�q�a���u��sUPk �--*����a�-����v���R��0PШUTթS��P&�+���4*��$w�=��H�0��%��P����$^�,;/��i�����|���lu����۶�U:~�N���
S�^���Gk�_.Ყ�G|�/�H\�E�
�O 3՛�" s,�iN�uN>,f���t�&��)ɣ�y�����-��5px���/������cSD��7&���d�\�1Q�G|҃,�A������"����s�:���6�j�<~���whr������HjvՅ� U���LT+T'�OÿK���9����2�c�{���1TR�A%��Jy*V�p7���8��tï���l}@eM{�3:e��L'�e~X�Gq�4JV`���j�q7![j�b�w�u�U��>�	�;	��E���cO�����	F�In�B��[F^�~d�?9�ܚ�/ee����=��%���8Ւoc^%�b����k{�x����˕s�pIC5�R�#*#�0�U�Eq-��������ƊҀ`�V@#��~�w�	�.r����a�թ����������jo�'��*7�f����C<�[X���:���( ����^�k۾Ț�ia��2m��Ⱦp�Nf��R����U8��Ҝ�+W��#8Z�I�*�
&�=5D����X�hN2�˪��X�F�{����xt6��� ���N���H嶛��k�ðf���V���$�	��'���3>�,� f�����c�S�Aڙw�b���72���ǽ��2li�<�s�+ʍ�N���a�Gg���>�pV��~UQ�����4<�]���5_���˔Q��Qk�+��<���2 �l���,'�򸵃�{����Ԏ�u֩4�	4�@�mo�g�B���/�����Y#�MJP�~\yA�SN�C�M	��~�%<[jO��$���-G���Σ��M�.��|�v������a6�[�C�W�J?��U���b[�>\BVu���F_�W`%k�'Y#9�I�p|J<^bé+�4\C���<�"��h*��Sq��w��^����ꨶĦ����9"\YX-���D��d+%V�)�.(9������v�8�d,6/��