XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����qȱ�T���< ^ ��c�d�����T?K��y�Ϙ=ɱ�-�{�0R��jLs=�aQo<t�]X�O�/v$!��/�#���ړ)�;y�&?�U'E�0V�`AI�䑔
Y�/��T����E�~��.�kԷ۟KS;�I"���h�j��}����d�tL�@k���#�YS�b���ʾ������R�kLs���<BO��q�����A�� �k^=VT-+�1�b��G���t�g�QP���MF�7d'SdqK�V-E�w* on_�p��8e��8�:,b����+;��;2�O�a���,��S�(��f�����k*D�9J���	���nU��7���mz|��$M�!�+�DKn���}�eo)�wC��LB�sM�멀�H(�Kw3韼��n6/
�mn�"�!�3{ӽ�;�Q��P#�T�Ҙ��T�R���J����{Q�B1̈́( +� ��6�_tgF��=`BKLh&���Jg��^�;r�!5�@@��)_޻����Dja�O��ev!y����no�"��d~��-Oa+#	tu� +m�>�*,�π�^�v'mv�F��@��)����]�~��J-MFQ��#��n�8(��%gț*�2���j�kh*:�\E�bA�cb\-a�vm�3�,�/��ȋ{����SZ�~ A��2ad.�\(�x�dң������ي�!�
?^bX�c���U��e}���i^Ti�ƹW+&�Ms,��o����9�����0#l��L�97S�vXlxVHYEB    2a4d     c10��F�V�����D䣲:3�>������@��?3}Y�&�����m"�q�6z�i��O�NK�!���4~��8)hl5��ޟ�m~�=,Г�k�=�4_�8�Jg��>9�\�<p��QH1�"�#3�	;�4DY��pZU-RD~����E�q�W�P���&̻Wu^d�P/��h��^2s��z��J����K���MtGe���ȃ���'$���/�HB�]q,q�co �RW��.�7 ��Pv3��X�{BVY��\4��{<�xX;u.��o\f�Ζ~ǐ�7
�����Q$������q��<���ax B�q� �s���3Ϥ'���[ŧ��4����S��8�r�G܋���R��'JП��R�t�R_���}SD|�f��Fb5�>Ed�R��_����7�m�6ӻT
Ǡ�ۙ�\ܞ��J@���c(�ʱ/�4�	W�J(qv*W��$'�_+N̄�:ϛ��1f��\���<����D���$&�<q=��N#y�Z���!>M�� ��6gӣ3�kŕ�8��׏ԭl�L�W�X�I�Z��k������ig��g
q�eIh4���a�Jc0�����){��u���a��Mg��?��Yej.w��"=�uZ`��\�"�zχK�"Vd	�bt��	*����@����J��Y�����1���
��$�����c�w���q6���0zV� $�GlaV$~�x�\�MD��S;�K�ItG��Q%N��{���`�@�5 ��SC޽�1&ŗ����� �N�?Zv�3�4&�4�oXEz�<�>e7D�N���J�g:�P."w� ��?���Z������	:��Wq擙<�&$�\>��|�t��k~�_�A�<Zb�򇰷��.9kK�AΆ�l�w�Y��cۑ��wh���@5�a�v{����n��לP6h�`�@��1��*S6�o�h�I�t�I<�,�cg>d>�����7��h-���C�8���yΠf\b��d�5_�O����Iĸ�&bf#j��#��3�~�7Qq��Uۂ<FR:��C#Ϥ��e���i� ��G!���ꝑ��1ژ9Q��m}ե��a�
��n]�,��}
rs���K�%��J&��4�d lQ�~�C�kS��&��� )���޹�	2���=�K˓;����������r�jr22
BB������Rm0�	.m���!�L \B��]%_�HL��R�QC��;���~V��t�A�y0���`/��7-Wd���6U�Z]~֕wDfdE8�*���==��< "�
1V01M���~��� �~�$�ri����n"��T䯈����1�ж��]�;fh������)Il�7n^ؼ��w����x��z�J�\a����e�L��'���r��v���l�a�mҝ
iW-�sY��_J��l,��__�hT-�xe��ٟ+��Č�=㯫9=Kz�O.L�UȓȨ?ޣ���]���$�Ȓ���š���롵�Uխaj�>�@�c�cr��آ;��lb���1���SaʛOsɖM��x�H!s�>}᠖L� ��H�]?��P�Դ)8��#SyJ2��7I�|D"����*�Z2z7�Gj�d'���:���S��V�SH�06�L���`&J�^Y&����3&^��-��.)�<UG	�}�C��!��������l����i�}mxג����,�a*p�}��JD߸��8r�Ϳ�Q����{����;�y�c
Ň8ؙ0�L���=V�"z�PٙH+\�Լ1ObZ�K��MMb	f�r����%�#/*�m�7�=����D��I�aui��������P����f��ҙެ��ky{��Z��-JZ!8F��V+�vvڴ�L+>4�'���R�}BW0L/q����ܧ,�3%+�vE�2�H��/�c�,�el�+��=��J�#�~��zl��.�־B�D+K)�)=�I;�����j����@���`>������6�l��|�EEu��ܨ��i����S
�W)��:Z��J8�z3�s�)M�����ūa�4�ds��g�V�^P�?�����w�mb0IUu��b�����([�� ���7�b$��9�>nPZ��⬤걕�,�� q:����fG��v�8�ەdz��R�&H�p>�^�M��ؼ|MF^�4�JA�O���Ă�oQUΌB�tg�m'7��!���#�V�U��f�k&���e�o��H�������=�1K �u�ɲ@��?�lU��;V��F�x ����p(�`��x�Oe���b1��!sҗN��A��ݮj?����k��V�c�ߥ .q�'��2w���'Jr��qX�����"���0��.O��xPj�N��L� i,�?���v�U��j�|`��%�?,I4�:��
Ll�@�a��S!��2�Md��ǈW���w�<� ��֢����pee���h����pw�ꞎ�Q'�#߼6%���v�WZ���\�f,Dء�Y/'�o��Vڭ�;�Y��7���F�Hc�Jl���1����٭�S�$�#��*b�������>
��,v���Fh�u.�����)�C�����C��:.jv�Tۥ,%R�i�^y��*G��j 4�S఺�'\��*�W,n�	i�d����^�>^�u�We��� ��KO��l_\��m-�|��>��%�?) ���:�e'DjA��A��E��~�G����:;��_a��ybUC�a�y�6x�r!o�3���Y�G7χ�w/�>0�V�:�q�A;�<�s� ���>�5��d��iR��2í�f��P�6�8j���B�A 9�
3�҈?�Z��0r���Dj+C/8��"pƊ��%��] e�
8aS�yE>W>ŷp�2e��Ar�F���	�=)�e�j����W�CJ��X5"�TJ�w�13��� Y._(�d�������2`�y��/E_��;��0�e��ؽ��K0_����_ș�#W��\�mH���G!{�6tl"r�Pe��R��ͣZ����-��F2