XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�8�B����H���'R'S�����%�]��� i��@�P�ot��~�k�']�Qe�)���Q�ૼ��<�~U�!�׊�b?�*�O<5��g�t8m�t0
9���Om�����E:$NDN�}�A�����g��p�4�|�
�P���LBurՑ��J��MCs+aܩG-v�ɱ7�O���m�'	ݦ��4�\iP(����=瑃K�C�X�i�f�֕��LF�(��X"��EK�H0� �z���pW����f�_cC��Vx�/_�H��F���;Vo&e}q	D:HMp�(�a�1��S��A�_�I��}z:��#L�鯙4�{iR)+3�ڞH���"���
i?�B��MZk�̲?�a��L��I>l�HT[eS �/Q�������ꊾBb��ɰ���MF��Y���S�MȚN�����?8��v4P4�2"a�3�аk�+W�KZ!��K�0dN���
��\�55����MQ�x�8B듇���
�~A	U{7	{�_��\e����\�L����<�K��w��O�L��xH(�	�,Uͽ��6$I�A�{�鵒-%/f��}��=�\'b������ e�=v�� έ|5��Ç����^ȾE�))
�{Z#���o~�y='�u��"��q�V���%���f}�D�P�j���gW�; 9L�x@�0���ڦ�[���1�Y]zkk����X ��7Ѝ_�?e�y����i��IG�>�":+��?B����H�!D�U���06Y����XlxVHYEB    2b39     b10������S�E��F����Cn����n<���H�$�
D>�3��7��8�U?�����2���M��@8Ɇx���Є�R����\5Y)�p�z�[���L'���TbT��[��� 3iT���_�,��y(mu�aǹ-��T��H�Ϩrwd�2!��5�]�eoE�su�ǆV�n3��w�"X�n���+>��Q�m���D*5]up�Cijp���o� N��r1��TF��e�7�%���W��!j*-p�
��h-��>��$��*o��š?�_���Fh���p,O��&ަM���٪nC��n�c�{$�L
�����5�P֚��B���Id�YB�nVv��c����>P�>�7���y3A�Q�b|ޤ�%!��aܳ�����t��U�z�r�j5��f0�cHA��[�	��e@�;�Q�T4����[���^m�(�y�}����w�ݣ�({qK�b���=�m�N�g�퉙.hĮm�#�\�B%J��=�����Gp���<�K̠�ʝ��a,4�[�4^	�*Cv��4�"vU��LI�4�@��8.�>��D��@��ŲZ�D��P �=�����*Q(&*U!�0�X�T��ڞ����TGd���\A�C�f�A�I���ηt#�����̽�G�,�e��H5t�H�x��{޹��]�tx�î���Mr:3Ѩ��gn΂ �I�8k9X0&~�Jv��)T`�?-��}��m֏�!m�B�Zќ��!0��*.#Q�T�I�� 2s��%�X5�K�������&�ގt"����L��C)���m"��j�?ᕁ��|�^ȡ�E'w�-�����g��,���;��g�Y���G>? G�x�纑X~��/3�6����=	�዆-U���������)2��*��ơ�:�
%�(����_��f�;��.t�������!�<l�ɩtt�w����K�VD��J�3��XT��{�jqH���EP���@¹��Hig}7��N��6��R�	�U�h���!���Ȟ����[�M�%K}�R���z$J���:ÚN�Z�R:�Q�p3<d�?T�rBX�\�9ϖ�b�T��NtȀF�ʆG9V�ɪ T��!��1î�����`�X���r��񖣽�dq��Ģ��	�ׅ(��H��L/-�x�xɊ/�z��=�
#2��zh�U��R�;�f ���"\�X�~x��c�w��T�}����� �U�m��(|@��-e��I��T*#p��~������?�����켴'��<hL�����&q��O�s��	i3Av&c���u�"�y)��bf����i��2g�P$�!�t�H�![�L���E���U�ns%+{;�E���w{���JO�
8u�dS�C��N�O�b{:�D�4k�Z4�VyN���4+bM�}懧�&��Cʗ�b8��ҜC?�H��R\��_�O^�O\��uN۴�]�v�sKбa� l� ��[Ӂ.�K;�;���zW��)�k$�9���yPO��U�	2�/`�l4��R�1W��9�+�{��C�6h)�/9<v.�� �<}=y��$5����[�.4���x_�oj�����i?i���H\��7s�&<+�Q��v6X��ӑDv�=:B�+ǲ��N��W�3���%}��,l?��*�$B*�����}ҷ�M�G�+0#z�y�H���w��d!��}���c���H$�%G^�Ǳ]{�h�,��&A�td@ap�p�Dvٙ�t���+6�}L�*6C��T� j̎��g�m�x�<TP���u��F���U�aG�%2o2)#˻DH�	\E�q��Q�1{���ۑ�[��L`��m�5�X{&���"�ǵ�Ոod�vB�%O�3^�m=�	�|����.�f��g�U�n8;&	����q�44Zv��MS���?���˨�
�A��s�7Y�6y�f�}�ڊ��j)*#�P��U����X⋖�A&���d29�m�M�4�a��~�B�� {h�W�k��,w������~���2:Ѝ�\d�x�Z�]���j�YQ�t�N0ۈ�R����oV2�֢7}nُ����������$%{�uѣ�o�l-� ��@1ѯnn�v!&��2�#�p'Q�.XYq�bJ�Im���i(J\U�k�T�:���8����#�T�7�6 (���jD�5;��9Z�����)���Nz��?�������������L�{��� w��}y�4��*M�M�Ig���(�9����u�M�041�k�3�nb.KbF�ْ�#�{r��3���z_���0�������'V_[�{��X����<en�2o��7XB9��
���,���څ����[���Liʴa�����(>���#�Րۄs�Q�.�v_��l�3��+w]���Ǯr
w�0����J�Vj�7~N]p�֒F��߀7��94Ӭ�����rq�Xyy��cqc 4��K�E^�j!���)��|����{I��Ëg�!�������̲{�H�����_&s�Pc�� �f,Vv�;����"��
� Y,��o���4X��\ŊB��2(�TԵE	&X��I[H$�%��T��X�ڎ�R�2u�]�Z�)�q�JZ�Y��.#w&�˚���;g�ӥmҏ,��w�}�����!w��d%��)�� �0��9��D���*X-Q�m'�ݝKp�a��I��U�O�����ɱ#�b������2�d�뚉p`9�T�Z��X!zUc�+jٗ2;�[?�P�^"��,�����\>�{P�ȥ�#a}k�{%