XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z:ϩC8�r9�fb ��7�K�6T>ϵ�9���#'�m�����(J"��҆Α�K�(Bt�^�n���I�5���9�9e$��[TK��z��
P�\|�-ԍ��������$_�Ig����?c{١���N9�0Og���ª4���q���S!a}KS祍��R�z��q���65��`\~2P�DF��4�˫�Y�j'�mV��o7�z�Y�  C]�{�8����rc��t�<����mT�z��B�d��W�/T4[��>�mxTgid�?�BXҟ��G�Gt����o�[�8��	_��)��h\��N3'�3�Ĝ�Vq~�b<�b����r|<3�9�F��h��n�x��v3?�u�3ka���ʥ��/'���#���6�EgfX�B���G��N\�X�#B`hg�����|�O��7�Nze�Gװ�Qr��R�hk^�]l
2*�Jmo1��y����GC#�?���(x}�#댜U �r�6���CM�"9�����C�T"%�`~݁tT�o����֙z�Ժ~����������ˣ:N6����_z&&y�;�,Vx�`X�d �V[G��h
�'d*R��s��r�b�� ����@�圁9�:������#	F�r)�Oo�$%�D�X{cN�Y���Ҫ�<�w@�F����&#�!�C���k'�י���7"v�UÄ��S�իZ{�k�C6��S�-"��#UK��%?I����~޿U(A�Pa|������ܽXlxVHYEB    33bd     c90�G�v���,!"E��A�}߀H���F�f[<P%�+�8Ғ��9��9w�24�a/r�fF��!���_�<���l����Z3(z�(&ۑŤ�V�-L�BVW3��]�����rN�R"Or��<�#R�����R��W�g��D�ꀐ:~�z�[ ��yDǁ�o3!<dw[<��7��s��N�^v<�ǎ<�N�����*u9EP5�0�z��E�|�|)�h�o�\f:��SPNcȝ�eQbc	�/N�v��H`�9�.� ���స�����@�Q'��8Z"M��ht�xaˎ�~�kɀϦ�**Kt���������i$"��1�δ��OJ~��i�(8�<�-�5���R��殤���ѷ����}~ˎJ
�:�hͥ�ս�7^��ϡRu�`�i ���V\5��4�;�k���c��"R}G7uYLKɓ��b��)-�r�7׺T��	S���=�W��e���k���a��F=�F |�I�;�[��n"������M&"��໏8����[�T�dΕ�ח5��i�����8���Q��*$@�X<Q�S��<Ea���1���w���z������l�I�#ޯrw< 0�Qu��ޮ+X5�o����5��(J�1����j��M��>�?�C/}^�`U�%a��y{����T�uE�*�YĘh_f��@G�IP�xJj���Mu�Q������� ����~}�H��,%I��=��,��~����B���w������� ���=��@�����DN���-���~RT���3A�V�e�/���j�uǺ
��	6��M�m�Kb�R�u����a�#=�[�|�n���n�n��.����s}v3DDW6<�	�7x�mt�5=\M���Ȕ�qu��M����� �8ڞ���0�|0+p�l�_����٥�y��T�����lkV�E��q��8�'���dh �!1�Ĕ����
���B,����_Ϡz�k�F{/�q�!̴bϡqp��*9E-���<�!?|��\j���^"t�MQwYq=�������P�����9���[}L~���9�H����s��ٹ�����2��~�p�o��ؘ��B��{�GO�#-��hcQf��oƚ��9W7����	N�nM;�������6z^ҡyG#7!��� &E
�	D��m�=	s2��� X�$u�-���%�僲Ջ''>oZ$n*tk��pw��s�󅇦�Hr/D�s��G��.D1����b<���?l�beӒݎL~�"��8�F���"_IJ9�+��"����^��HƵ|s�0�����v�T�m%�9��/b�L�p�ϣ���������S���z'�M_���f���1+���J�+з����|�y��ԫR��[�R���t;K��2�y'J���x�i2�l��O����Jn�8q{>Y�g��J�~���1��f���V��)�]�X�����"B����v�Ϻ�O) rW�\^S��fDB�/�)�T�ƃ���<V�0���݊��+�/,8�~fz&f=�<Ӌ�V����'a�	O���_���Q���a��J��~t&լ���C���7��r���z=,H�q�<���@�m�RL�㌦Z���ۤ�AJ"*ڑ`xH�u�=�9���<| q�����֭���ٗu�~���zq7N�Q����jB���T�P5��ϥb�}�A��/��k�(�sWΔOQ
k��Y�Oh�ȼ9�[M�V!��3=6�q|t,�$m�a8m��K6;�ms�e��u��r�wx����BY #����w�W���v Fˌ;�� ?T��x�ߌ%g�J�Pr `rΰ���x�ͤ���s�7D������0�2�B�m�QY��>x��ʄ/��O�Z �^ѧ��d�j�X���O;�ũd��'�NV��H`b���i���A�h�+I��nhx@���Q���J��b�4F�9|)`7� �n�1q��'=���S��x�0K�����ʒ������P�$��S�x�O>N��o��܏��r:Х�ظ�E�0ޔMw�c�Q��9@z�=�d�O��|H�F�����j���4��eQ1��Vj�F�:����Z����g��n��8�����'ǒ���5�&>�x��|�]�C�9l^�\˺"J����-S��aI��'k^ {����ۿ\��s�[��2�h�+۲[8��#�0ע�}rN3K]�:9c����9HA� ��B���Š�s�V�<�`R�O4w V��8�`�Xd����������T���D�,��<ZE�2(r�����Tr��0���ׄ^��[�Ʒ�9R��Q���q��8�Hy������{�o�&���]���l��xD d:�ɒ�}Ǹ���?ZGX�Ѝ�Y�m��u9�u�Z��7���}B���Th������~݃��+H�=?���1p<�x�3C�{�N2$���<���M��z���[�0���HW��rޯy%�9v���f(&�8 %]f� ITg�lv6��uu��/ł��^d@��`8Rހ�_!$�YႃVQU�����ɺ�8;R�N1h�z�(�+���s�B�k%�ߺ�<��I�X�����!��F��V'bs�Q-W���;?!�a�j�����6��O��^�$4:fI�P����:�ı|w���Tc3����6Y`�a�i� ��1ķ����Fǩ����H����ݖ@����*;O��$��Z^�����/�J�Y��y��;_�r��0�j��:݂�2��/�8k��xG��
��z����4��Ux0�<g�;K�AN����a�!�Q�Gh��izr�^B���^�_������\OE6��)��Z�b,�/6���`�ӝ�*����/���?�X��3L�����m
�_jl�T��U���w���O�����^��J��,�cmj�=ȼx��j�\�&� p����o��mϚ�I\�󜖐K�mN�T���@^�U�%.�K�kgmJ~��#IW&�)ݽ�}���/���/߽V4緮L�!:	��}6`���kai�y�ȈvT��9aZZ�w��2�_����r�IH{YA�	�����|;=��6a�5���/��ST��1��JU��E�<ۀ-,�=f����I܉H$`+[-�%�7-��ē��X�j)��b