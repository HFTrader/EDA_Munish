XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8���EY�(���X�L�Ј�n�)C �۝Y��*3R��c����g��Δ�x���S9
J��9��Z�K�޺w�Ao����z�� �xh��}ޗK�L��k����X��B�<l��D�>ˠ4�4�=фk�bm3��Z��J�I	��N��V��TM��a1�^�j�9�1�����}C�$��� 
L�H3 7=҄<�#�L2�3�wYA�!�lH�Z��E�̅_�ţ����VV��z��\��[�=]*�%K.̽e����5w��18]e�"�z����{�<�@^*�C)�_30W䐟�c�{�r��������Ի��
p�o%�WФeL����2rI�%�:����6�$pl��o�""d��T�E����N+�h)P]v�82�d<���F
� �O�뿑�d)2L2a����P M�f0������%�1TT9:򂈙 �΅z�/�(��r���?J��PT�(4�;{_{9e�q�f�ۀ��J���$N�{�^��UPd:md5��bbsT�u[Ԇ���p�E���V=>�M�Q�\��d+�kŵ<�C� ��˱KT6k�i��,�&x�O`��Q[�ɋgvl�	ʩcu^���)ȡ���I�����7J�Ea��� ���6A�� ��{fgbU��<[��F�@1LY��)p���/����f$���ʆ��W}�k���.���~�I���uQ8�+�fTO�묝dl�7�|Ci+>�37x2�#�!P��W3�XlxVHYEB    fa00    1790D�����n��QZ�H�����6�b80��B۟b]�nh��ST��A2w��e����DH�C�`�og���0�7�sW	Ɔ�UT �ǧ�����7P�\�-�!5�C���;E���P�_��x��g�]�v����b'E��k��ߞ�	�� �a�G����4�d:�`�.����Y�����)�T��*'�.�tFÚ,6�u�
D�O��JJ�P�U�d�3n��Ҕm[���I^��1ǐO�5V�
-�[��C(2^^m�^1�J'���[����tߙ���Dbe?��}T����|T���xs��Ec?<��Ԝ�7pu�������.7�P�D�:��m6)u3���6��iSK윗��Lv�]���L�^ ��~v��'��Z�i�Y���=Y��ֵ%��l;�7�����+���XS�R�^cr��`��#�q*���$�b�b4����"$I�;j�8��݂�q�=,g ���č��{@Z_$�ہV3@����R�L��S�DacK�|�p����$�q\jq�L�S`4��\�>�U1C�$�ǁS��f�a^�g-��C�;�4�[��D|�o�'ܝ���Ř�6��ϊ���-��d�z}ƙH�>'lx���|�� ��"��9� �}{(���N�7����z�Bk%5또2��[Wlx|�����$ �#��l{M�q�>9��9}&֟wv��q&u�m���Ʊi~��ucxfó�/�|���W���b��h��xr#�=�d?ȿu�����7t>a�ԚY���Ese��A�w����k���p��S���l�.�4_dQ`:�/��WI�H�R5P5{�ӑ��Us�'��d9e.�BS���ԧ�rO�h��� q�0#$�&s��a|"�S��ٛ�����E�(��D�?��i���'1�ɟ�/D�J&*�	�'���Ql�V ���0�±T����[y��*�\T�d1n8��L�h�n�	�s���̊�0z��\���w���}�O�t8��D�De�8p�ju�̞��|���<�I�D��&$2}
�6�z��G'��adj�+cz���aĸ^�3/n	v k_���F��pa�=��7C�R���7����?��D�� ���{��:쭇��K��yi|y���R���EP��l� =��Z�	��i���y�"�I���b�a��?RU�Y��
���M��>d����qs��NE9n��wmoSo(D
Rwm	AjP�lX��������Է��C������ٱ��H�N����/t����ˮ	uZo�����^���1�����e��S?Ҵ�}Շ_O��D	�oN�[��KwU�
9���	0��9D��It�;�xHc��.Zi�7I@���/�Zij�O��G�L�1`����?�w�/p�
[$�k�ψ�;����b-"Tߘg��{<�DoS��S�h��&�&�Q�O8�)�%%_���?�k��g�n0H��
GS�����| ���m�K^R�	������.M鼭`�?mHl]������M�u��g�|���u�y����҆��a�Q�z�?���F[�J_ԯ�]�+.Hʓ�����I�#J��^>p���(��:�����S��d$k����V\� "y�"��3"��gM�Wқ[x;HwS�IېjT�;���SX��y�Gc_=&ö��]�r/	�`�����{Q�]C��ε�;���|:�� ~3Z�5��R�q1ؼu�L�)�9l�%�i�E?������Ɋ��� @����l}�[^ĉ'���R�x�3����~q�G�|��hj�f�|�;(�fǽ�3��<��r�|���������2
�� 0��ے����e�F+`���t|G�AK�t�B�Ck��هH�)�,�j���H\��N��|�%��8�A6��D?�����׆��M��{4��%�q��6ښV�k��}p����$q��n�p\F���Y�g@���ߛ:�12 FVu�6�؇�LJ[�^??�Dգ�[�y�>,qjy��܌���;#ɔ ��;���C_k?��8i�M:�jh�uxg�7�v��.�@t�����]Z�,�D*lݻ��r�R>��\����I<�	�r1�V-0��`�Umj���W
W����X���.�4h�&�3��� Ŕ�N �� ���/�,�̢��C�&��l����̋��~�
�v�3UFzC�32�b�as���!B�$�~ �A�ܩ����yWװb6�IH��En�@�oF�:�+z���'�~�����e>�_�99?ݳ2�C2"η_F;/pY~��6�є ����xT���-���K��9���g����aܤ�f��04z��*�N^��x�V�&�:�h�&��9���`�VŁ=���&�{A0��k6�|0y�!v2�H׆����^$�ت�/ڃ,8��Ĉ���cÅl�Jf/Mb��N��[�=n�)����Z�=�����2��ʽ]K*���O��g��ݐ)�{e�'�~kXO��O��/cvc rPg�'�8;��{^��SX����(�����5��<=�����-4�6�J�{PF�?Ac�E�0X܅���������<�c�y��-����[�*��;�3�r=e?:E�'%��`#��A���%�����s:@�<�^�=kv�O4ERUG�z��)�y)bRP��}�M<C1��zױ�:�%��
6`(�R,��$�Vdy��Z-����Ǚ�A��<UF���֤���
��	g����Nߦ?+��r��^>�&#��.Wn�w�� Y�@��,�i��=U{��z������rR�nӢ/�;��A6U�7.�����U�T�$�H�rV��@iX�_f�@R� R�T��7�9���۫{��o�&�U���bD�u���n�� Ѧ�I��s�a�S������U���;�3S�J�W��Q  ]B�6UGA�=:&5Jv"�"<���g�驹�߷Z3�hX5�)������м d�������`� P0��[dL�ʗ�U^�~�EfL�@�c�N]8��&1|#��p:�`T�^W.E��p~LN&Nt���h#x��c��!�#��,��
'7���C2��^�2���;*�`Э��!�k�B	-t�U�nwn����O$zFT�)�����T�
݌��
i3��-��f�=��3����I^2ss��`��#α�Oml��V����R˄��^}�C���~is7Tʸ)K��.�6�Gt�K;��	o�1v����[���o��0�i��Ш��2o}{3�\����IvA�q�= �������I�J?�����Q�m�%�T�����&k����5/H�;�f�-!ikvq2���I�@M�LGCYȢ���\��\�`�F�ci�Q�Z������Ũ��
!'9�R����������4 ���j�m@+H�0�l��ƣx���}��8���{�L�1��{���'2���/�&�-��/��P���D�(aFD�j�f��E��S�M{��V�r$ꈺ�r�O�6��������|�V��l�h�����i�1�	���ї�wΉ?��ũ��d�(w��_p�]�\<,!㞛�v�	El2�$�K�qv�J���
2�0ṕ�&�;�G��x4ԯ�]R�a��j��N+t�C2���K�By�s�m�hx�-0R��)���`�}@�&�+�t���\��P��)� N�CͱRlHp{Ē�4��F�4�x��/4M��ұ3� �j'z��z�bxKwI��w�)&�B��P��<��5�y�r
�Ð~��R�0RfB p�$�4����Q~ ���9@N���1����7'�*R����[Ɉ��9��Ӕ�U�W�}��7]��o���鋞�`q��נghOf㐲5!������ۍc!�Ok��rw=a�9yq���d��y���z'e,{JX�
�:���K��Uӌ<$X_,���`�������T �]���и�4��΂�	ʗz��G��#�l�c����N�����4y�a˶{�J�8����R��6���?݆ǯ��"<�L��R��)+��?Ƽo�Wg��^��{�������6��z��i���~s��K����T�Q�5��Yc7h.,�����K��ZFB3�"��,ѻbȘߞT����y�o��P`A�����1����jK��p�o-��[���:�g+4�y@0��!�u ��Kec3Үl�V������{АԜp�j�t6Ob���C�]`n7Vy�M��0����-|�YQ�9�V���1v��m��=O�ߧ���~�2�	��.�g�N�E#%;m1�n:���.����<�__?�����S�i
"�KG.:�4�IJ9�U'���F����lT
dڳ��䴿�YǛ������Nf��W6_.G����k��|g�z�Z7����9<�'	�7E���L;�X�t��~��p���!��l5��t�j����"w��Л��v�ِL?�U�W={��"-�J�0i��C۱�*D_��N�F�>y�9�b�!B��T���gp��/uw6A"a�0_;��x`rgx���������!��`PM�o�?:��`��%��(�!�|^}�w���,�F��u�S��PR����a:��Dv[p���� �IT����ciNٿEGr�`�5���q罙)� p�u��m�@2�u[,Jʠ�
�搽΄Εs*�3Q|*�0K�3���W�3l_P-/מ�$����!��e��mb�9��"}�2p�.��h���AW�$#41�q�>���s�	��n��v9��f&���|rU��ԇBd�]�������<	�`�Sշ��e`76���,#�d�&m�//��^f}M���u̾�j�q�V����0���>��`x,P�`%�t��v���N)P���+/;=��^�iRm`UG@��%���\B���+��l���D�Z:+��n��e�j�<��ATZ���hl�a����> ���?��٦Ci^�R$��C��]!�p�eT�֖�!����21���Q��?��yKj^!������u/D��>dY�ZFI	7�m���5�F0��G�Z��A(K}���\8�G孫���(0���a�86YT�}A�Ρu�\"4�w���%6��Ӵ�z��͝<���)|L�۴(��e���l�g]J}����|;=:6 ��)���H��,/t4V}��)Z�V���(�R�!2ĝ�y[�n$gf��k�@��@��֧���V\��J������$�,����md��3j΃#��9�ؼVc����2�M2c�b���i����e�#N�����K����g����$�ލ$+����,lٕ��aC�y;�*ZМ�HE0pH�z�	*�RJ���� ��$�At��+��+�2�\Oj.y�J7�gy.��i���]�;�9-��x��#@LM�?�;�&����W\}�'%��&�����c,�W��6".P�������n���-����ά�_�z=�'�Vr�u�sLa�W�dm��?Xg���LD�ɢ�85*]Ӫ�~n�"M��A�����c�j
g֡MC��dBΔ���|u����eJR���^|�\"�c�g�j�,k��9"�?���?���pe����T�r'yA����b��jE�+�����;!����_�Lm�Qp
�A���t��H������b�zڒ��[1d�ʖ%���Y��Cޯ##�C�Q��]i���~�Y�'ɣ�;�X�ĕ�}�`�3ô�D���넟���0գQy�dn��	�H6E�0��l�;l���}Ӭ�gu��_��v-����FN�i����u6DV��_H_�-����v�]�0ף��xl ����%*�YiNk�ϙ8啧ݜ�9��I	1�ù����vG����>�l�sH���u񦆙$9]�C��6��.����XlxVHYEB    fa00     5d0MVGLdsQ�yO���Y�!W��Ks�#��ڷ_5sr&y8���H zq؉"�3����(l�ۭ��:EI�Q3ٷ{�SPK��|�� A�"@�i�gi��U��qF�/�k�5��{P���Xj�LΠ���X�`�Y )]����h���?�-���z��3����o�F��f�6=8���q}�$ �m�0�w>�!�%�V2�6_�u(ѝ��<�����xY���AlWǐ>`��woe�sٜ Ӓ�F���� Ƿxz����xy/\��i���c���tFD�U���x�FYf�����D���c��m4�YU2��	r��M��ީ��՛��\6s�����%��΃�����BXY�A��d#��ʎ�@@(��^x�X+`��B#[���z��l�)Mkrm.L�y�Kި`��B^�����r���Z��O�3q��e��,���>w����d�i���S�[�m��<P���x��kMq���j,�RQ���xv��u�V%�n��� ��!|G�����R��t�U4�8S�QCbWC?ٞ{'A�Ϭ1�����U��S�;����F̠k��u�\X�DL���v�!u�?0¨"�Vy�c9��ͫVk)���Y����{��vV��T�q�&�X��Ռ�@��5.9GiPĴ?��)���5[�qC	1��bG3�0g���p:.���i)��i=r���#
�ZALD�<Vsr��s
�K1=z�̎7��Te(��%$.*����柆 ��	7@⹲M�l���Mua�Wy
��u��b|�����	,�'^�^���� c��f�@y�C�i�c����A܈�7Em!�<�h,�x�EBD�引�K'ꠖǞ3�O�»�d�r�s7��p7�
ķ�柁�
�F�^�{%D�Ü�k�{N�\,@��zN����mĨ2v��ȍ��}�U�g�����Tly�2�-�r�;[���h-GzCÜ�����0�`tgpi���{~���o>n&T�(9r�����=�2R/U@�� �I�ų���ƶ��щ����� �+�v�VS�P��7�A�)n����wUy#��10��O�uE��[~���G��䢍�ڧG�����Z�w��.��l��L@�n7��yfBv5�m��߻f��L z���t-���#Υ��^ѷb��c6���KYH������b�AC�b�Aw�eQx���f�$yB���,t���5[z�g�)�b�����3�`.�����f��+Ks�׻7v��JBYJ�E�9�Ŀ�t��R���r��[�#�.�b8($����)�f�.& �ܙ�<&^g��~����~Y0L`2��W�L�g�=��Qpy.����<n��8�xT��B��́2$J ��VhM/l�������k�6,\�̢lw�/1h|E�κ�u� ��a�����5`��ވ��.�a�U����|���2�/B	sS���f��v$ЌXlxVHYEB    fa00     640�K|,�l����N7�x�N��B8W�oai�j|xX�Ƣ{P?�=b�,U,G��F����|ָ*NU��rh��ͥZ�-�5a��G�g17�u�,�H\X#���A9���s8{~��r K[ٖb�z�����|k��u׸N��'.�1#y��]����9��a��)Y�AI�;�?�'*%�kyo?-��.��'�%�~a�О�*��;�	�o#n5L[z���Yl���\�!8fW�����ǌ�֕�QdgEt'�"�'$p�m�I:,<�!_�	epӹ���]"��c��jw�ml��7ZS��s6=�������6l�^c4H��xhRU?L-�u{*?sr�,tKϷY�$���y�}��'k���s�!��0� ����_re��߶��F��s.S��X:$u�ʻ���]]�ԉ��J#^��Xg�[E�x-�,"ݜ�vkZ�Cbo�ڞ��<&g�������Z���3d�B�Q�ٿ_	cn�W������M����H���������
���r��LQܜ�����h��'>L�_!�5cm��C�
�x�����p`�����|�鐙��#(8�d��@�ƚ����O�NI��)��]0�u�{�ay��F��Po@B�2��x8�$�\��K"��ø��^�ʹ��9�ܝ�Z@�p'��"�2��6�\��������lU�����z����B����������Ŷk 2����T4�$+��R��U���|�C$�kQ����6~,�H����H�/(�u�BLy����.���:疯M�WfIL`2����vY9�:iY��H�J��Z�w���|"|U�-%����4�V�&�^�-'��G>x΍�)�YK`+�i􃳣Ʃ{��G8	~��`a�h!��@�d�����#�3m�tb�R��,�����愲�J������{lc.�$���M(z0J7��P�zM�HP�e"ϐD<��7�Y�Ne�w���@
��Ŋ�º�}��5����L\x�Z5 T��	U�7����G#o��8��G����y�گ]Fj^|�����j�8�1
��ÃS��";�'�@byƧV�SH?g�!���,����@�7a�96T��?��3�}�n�B?��V����`��3#��jⴶ�ͫ�`ɜu��ɗ���[�lIT6��)��;z�cp�*?�3��a������;�n��c�F�
]���������zE�v�qVoD���lN�He:л�	�o.�)9�Ń�q��%8@�����P�bw�ȕG�O�9i ۪�(5��#?l�w��@c1�"��v��a�:;/��V�,��צ<�A� �=	��G�w�i�Ҍ�}�<���e�Ԁ�0РAϗD���D�Ն��#��QCv�"�|��AO�:�E'l�x18/2��?j�}���Ӳ��b������t�Y=����]0/"�y�06�\S�9��BTB=��{��6H�� *WT�����_�#U�����o �o4`F0��S?r�΍�:2I3��.���������l�,�  ��El���ɝ���Ϣ�a��h�e������wѮ�gڰ���A��}�
���-��狍XlxVHYEB    fa00     5c0��.�����ܜ���!o���"}��[Y����g�����^ܤ��ē&��أ�W5��\L�4��=�)�!�uhv¸�tld�EY�0M�Pc5|n�PG�(`m\ٚ���֘4)��|���f�^�3^k�6����k!��	��X��/Έ��	V�Ϡh����CMA���J���L.D�|�p��AX(����x<t3Q)ŹG2|�1޺K��,�ggG,�e�cP���ʗ��Dͮ��>~M%AiF7�^&��ې��$��X����r�%�U����"�x:�ٳC���)�XqЃ�cW��͇o��)�5IcQ����G��0�Eҽ�L~�m��8�N�i|Q��S�
�p�R�[˪�ka�w�.��Tܦ`7�n��5'�������D��1Ȗ�oؕHj?��?�����_�����7Znz��6����3�#�勘L���n�O�Bt?����h3Ō��,�&F��D�5+�VB0�� z���E�����`/}���˴�׈��򁼼jH�ْ��*���~�/�MWK�<���e[�� ��I�EaK� �`�c��=�����8u������ه���~�䓔J�7xjC�2yN�2��Kc��]�:�e��iܒ�f7Y��vWMo��e�� �e���s�:"��Ku�8l���:޾̌����g�*���k�$���J�fdj��$
�6��;�۝���n�ޱ����L�Cy;�<2x��wJ���
�F��$6^Є�����ah�Idw,���rMK��� ��L�TH�5�nV������� ��QZ-�$\E��[����+�l茏������v�W��	_�0+ Pr1F�m���91�����-�@����YO��pZX�f��?Y��>���$��g��ִE�Ja8�2�V蘔}:��n��}-�B���� _���Hae�m(�Qn�:�O��!�j��0*q���5��d�y�P�E�n]*_S2�U����� 5��!o$�&� �V�/q�8��X��z���P�x�c��aoE`��9ڙժ巂�Zx���'I��~���#,UCF�xE=IV�5��Mk�)z�ͷ�Y�6�%�X��3wK��|Μ�z胑�s�b�r(U��E�l�;�+Q�"�7m�ٮ��&��(��0�/M�N��sb�ob���۴�s���y�:Ʉ�J`='r����&o*o����i����������u��<�u�s�8?�NA�U[�	Y	�OU�!���]���{�v���!�fX0��/"��j�Y��ox8y|b+�[���O�&�p��LQ�S�m=��{u@>(\n\�o&~Q��L`ߐ�����2�ʲt4��C�H����ch�B;J�SĴ� �x��"(3<�XygN��1�$i�x@d1p·tCo)��e ��t*�x���۞�z����^�a6c/��nx�C�։�|x�XlxVHYEB    d347     a90��j�i�� 	љQ�5ǮKX�ĳ�tD�����iY!$M:9�
�ԏK�����;r�Gӊ�HRXY/v�]5�Ťf�tD}h������v�WT:��[�}~;�X>��}�'�dne�8#�gD�6�0ğ�;�r#rX�<EOf<jQ7��U?�#�w��Mm�U���:�<k��@%W)��V%�by5�kA(��j��[`�_˫Z�/O��%�=#C@³xnӼ�)�zѤ��i����3�y؋ص��� 3��Ǖ ��C�J`�_��ĳ���Ӣ���#�d��׷�*���n���X��]�}�$Qe��^*��ֵ�w���̻?U�WU�r��ز��-Ճ�}�!��j����`Α"@�ke��M ����y6���Q«��%mM+����.6�6վ�B,��#���\4k�k�͖��&+M��n��k(��}��p1�b=�*R�1K�`"b���w��A+8*|7. �bP;`����PY&�V/p��}��WR!o �O����hЌo@PL3����VaFG"@��r�(<ـ�8
����F)'��9�/�p)����i4�Z�j$��ʵ\X�����$�[\TnA�#]����E�Sع��Oi�=	�if�;�ޥ���,�Q����%MPGS@C=���a'���W�:�Q�so�}�؋P���v��CQM=�la�ME�e������XE��ڬ�r�����_#��Cu8`��;E�"��]�X��dC���-%��"	�G�	M��Xw�D���")�j��l�����������?+fޫȺ�ۗ�:5�Z�|P�2��[57� �2�R�
���P��Zj���D��^���B�$�b���֑�y�â���ZϽ��L�Nw�� �OPq�?�ZI�cԛ�����������*�#V�VN��V�e�ap�Y3`@�Q(�!tԏq[az�V��h�3�<�1nT�����0/�=�P�xiM���	;=B�r���B�&�� Ld�D�\�I
�i�}W� ՜����@��=�fP�zHxf@𶣧&2|=��<�+�!)����8_��<l�O��,:�w�Y�<_!�������<�[�tF���h$��V`�Iְ�0A��P�o7��ra'�j/� ޣ�H/0:�Q�A���יQ4���K��ㆇa9����דeN��L��q`�,��}���ֲ����\�u�%.�oX��gF8��g+Ҟ�vge�`�p$���� �-	}���<�ub)��zB�:dB��5f6�}��С�<�1�sW��՝�sp�lq=��K=�w U���d�O`�S<\��@>�����~��]��kSRL>�$:�A���K�׎ϏVO@��d�W��8hi�5SV�����c�!��Z?��o�]�X{��Aj��o�Q�`		OK7U(vu!'�H6k����������B���n�4�������,g+�e���m��]�	?����=��@* ��}�K�UfE@�j�;'aV������Cc�>���Iȼ� ����w�U�^nF,��Ҏ���vcu=�I��'���Ņ&�!��eB����y����0�Ù�5��v>:�� ��N�IZ�K��A�z��j�QS�����3��I�� ��u�l�o=_~Ѷ8�(��L��.�Z��:^(����_��R�d6sI�k����+ѵ�+x$���蛢���"�@�9�/��Y\[����P��X��Q�\�q�I5D�Kf*�fᇄ�,�]a���`BsY	l��"����A�d]���}���P"D��map��_�p�y�hj��_Eͬ���WU釱�h:O%���L<340G�az�R�M[�6�r��>R,^���~'�:�J9��eY�T�y�"�j�<�cCɋ0�Q.���W9.��"�y���5�O���S���A�_^�ȣ���S6�؂�h���+�АANQ���	��]����V�xȄ���ft*�Ae��e���(���)��z�h�\��ӗ�n��k�
�	|�N����Y�g,Vԓ��y ���Z?��|ٟ�(;G� o�4�:�nW�Σ�M<���4�YEە�dv��F���C��^��3�Z����Þ��uC�9��s���LT�jo{�����t�6p9x(
�����VT�::u��O�^8򧜫��d��Fl'�/����r�<蚚���^�˻���V�(%ӕY�bO<��T'k�x�FD)�0r�UH`����FK��VN�l���d���V;)ã�X{��'�M�{�c(b��ٷK���a��;��z��b��Y�U�T�1���/�R}�V�zC'�
�l:`���UQ�6Q3(���Y�JZ{m�P������R���+M�u]��VBB��M�%���2�.�
�-
�����v'X���;���;ks*�.&���+.�?O�K���l��� �����E�,kԔ���T-�	�p5�����$\�yR	�c�O;���&�O��O�&IG6%z�A��/�'��K����`�B',�|PoSD�(�@����rY��)x�,uLlS�ey\݊\M�w�ȬS�˅/��:�Z��@��HgRW=_����z����j�^�*�w_��Bfpb�~$}�?�f��c�l�E���59z�5D�1�mJh�5?���=�  ��!~�5Y��������