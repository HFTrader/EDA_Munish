XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �Y~�h��r�J�c~��x�k���'�^�a�6&�=K[�4����ы�;�}cD>Z	��+m_ؽ��.X]�9�l�z��"p�����m��̉��[ �S�����2R��e�� /���Xb:��$C�Ї�ȶk��Q$�a�$�HǓ�Z?���'8q ���B��|r�<�a�NpRV�W��^C�J+�(t(����H����j�0�N�)<zu�m�^�.ßMn�"����
�:��C����M�Q;�D�����<�B��2����sp�-���Ĕ ����˙��	�r}lADweTR���rX���_ӎ
�{	��5��%g���}�FK�t��c�����c�O�\�M� ��=������6�x�@�p?t��FP@�2������֑X���?��4N�z���8��z�YW^bh���n\Q�H���}�t�#>���[�9Y;�eW'��8���0i� ��GjP��5AC|�F�+�NL�Qɳ��ơ(a)�&�4a߼��i�{�ͤ�	��X���b�+�_%&�a/�kP��4���ƒ���@��b��>��ZM/��6�1�L�v����6���]hn��#w�ʌ��Z��
���Ltq�Yu3��_*g�4�)ෙASrzU�/7Bdz�v�k�S����H+�ᘏ�	���%e:�U.lΣ��\���N��p�+�9�ߩJ�6���!��~E7��*y�AW�1����1�-������������dP2}��bχ�F�8QX��
-XlxVHYEB    6417    1280Bņl�"�<���t��2Foঐ3ߌ���<��R�Fm˞	�ͧY��GΩ���N�F�x��QO��-Sȕ{΋�t�O!:���!��~ґ~9�x-���snn����Q2Y������>fSE���a]Q�L��k��aY�����=���(��n�:bl߇�\��g�����(\��i�l���$.�hQ�e���l���>"�cBr�ٙϿ�b���j	gj���=sLjf|�x8D/�n��d�`g���'Ë���� ���w�z�q�Ъ����1Z�4ԥ�������$�C�`]�*ʀnx�Rs�Y�#�F���f
c�$k�'b>�m"�T^�%ȚQ��D�����`隢.T�3u�u���G�r����������hV��Y��^Q�dJ���Pp�t ��d�L(~BYڐ+���W3hط߻0��1�E�P�7��ۋM��
N���բ|�tx5� v�]:�$�נ�=������ �EG��y%4?<�8������b|�||�������3|Ж)�eʲ�	���Ed�v����s�!"f�`�4$��n�T�S�X���[x��M�yh
L�3�LE?�����Ⱦ�[8��[�hy@V��#;��L׊=���$ʁb����%��"���qᗱ�$wh�9ʈ0��N�y���EZ��L��k~&B��r����3�m5����F;'3r���?j���	���������f��KbF!����ٴv�|~��W��3��w�'s���s�#L͎�-���D��>��Ɲ�"�(X�^�I��J.zV�Sg���Á)����Ga�R�:�ja�S�FF[�*�N���k �q$}�?g��}!Q�N�B�p�M֤ ,�ho�
�H�s�.8;�4IM�L-��ukM���ۑ:'���f�������ˬ�N�D�jr�vR@/�s�OP����ز������˾-	k5jj�U�z��L�햙;�5�P�4��p�D�Мn~B���)��,5x{��):��ft��?��<�����.�Z��z����X����������Q|C�Y�ޤ�ujˢ�v��X��#�y|~X9t�B���6��[(�$���=8p� r�(4l�\����qEm�I��2MH���$q�<��M�B>\������>&�J"�Po�x�?/�m64k����n�YykJ����2�T�sR�T¹'%i���7}@*ẕ�5�����_o
g�\��A..8+;�:m�σ���ʵ����~îQ}o�s@��w3��T�Q��К���k1�]vĲ�Li"ĶCЅK�r1��Z(?���9D df����x�cH����2��|
���l�z7���ʴ_8��\8��̾ŏ� �iX+�������Y_,^?f��G�^�\�(��laV#E��6���ތ}�KV+�m��0��4a�	��-��/����Ɋ��݂*�J2]��y#��8Qy�q��z��?�{��'\F%�V����}[A-�ְ��4t�ӱ[��[��؂LVRX$]�|w+���x�CӟS�a!U����Y�}�_�1���To�>JM�&������V��[�l�n��wH0{��yN"�??&S3�h�	��3�ξj����u�J�����"IDv��A��/��L�$��t]��9�ۧj�!;U#��:A���Qi��A@���܌rj3T����;��䨽w&q������,綡��sXb�N=|8T2�V��u\�~:W��c���MQ�b�������>HwI����%E�"+pQ�HX����i4�7<��͓{���ټNl�6Ew��5��M���Y!����SW����vY�kK��E�!,N~�V��l��#OQ��MS[�-��G�3�VxV�D���y�S�Cƍ��'i{ �Zq.�A�I�G�d����wr���Dkv&c� ��M3TNJ~�� w���~�� �_�;�ur�^�!����{�`����W��v��������z4xd�x�8�ˆu�����!���'M4Lh��]�M)�����&�T�$8��{�K>�9m�%BA����Ӿ���ݍ�%q4/��h������½�>��@\��s�#ZO�#$���BUW�a�;;�o�R�R?�!J�AWdhѝF�Hi�5\���p�N�39�qfSk84?q B�e���'ŧ�Ԫ����JQ��ڙJ�!Ip�gHul��+��Qԝp���"@�M��Ǩ� |�LS��=���*iw�1�e�xi�������#d �XҚgn���g�K[���Q�RB'^�-����1�/��u�
Bѧ/�ȷ�E7[Ë����-�4Rb��>�g��F9� Ԑ'�V�0+��,�/��b���qncFv{��B&����1�H	
�Xi���IcV�f(���e����B�p�r,⑙��ԡ%a��U�!
'u�����;�F_�rd߭S�a6do�BKh,�~�i�|Ex�>`FS[��p5�|��������j�]{�~��􃋙����hN�_M.ߖ�^����K�GN���j�ln ��?�c�.)N/�x&�{\x�H���ʌ�c�����ֽP�p����0�Ť�H���2K���F�!�Nܴc=�PN��ǈ�>��
m�Z]��{8�Q�}���ת�?��1O��N�D�������G�
	�"���^���d�
%oM��NP�������'U�c�p�OO�7iQ�(�4���\�k��1�۵(�)�e_)�{�!��"�$�6tc��v��y�j����K6�w_p��q]��\R���L@�:Ww�F�Ql��MU}o2�
0�|���
j��$�Y���S���a�:=�,Lr�ɔJ�c�����,��H��cUX���ώB8�e��"X9_ =)��tO����l���+W���@����1�sy?m�){�������.���A��d����<����n�nIS�-M9߮b�ў5e@r|�w�T�z3F��Gs�q5��+�]�Yh�`*��+ɼ��)��Z�&���Ԛ�y���Zq��={����mPn���U����T�]*P�̯S�l��rC��b�w��Tڽ�q���T�`����M���L!�z[b*�~�0��u�I�Ǭg�����>$�9�ꮲN�w��� �Zn	?�8JuQ>J��%C��Ib��>��_+i$��� 8�G��� Q�������= �q�g�����s,�H�г��p�P��O�c؏�N���:�z�x~�*�*h�� 	��PC���:��6 ����ڌ4�-��>ŹG=,����K���)zB�?�����ڲ�4�Q|�	��,�s���,�+9��	��'�mo?ߢ�-�F=�񄴦l����uw������o ;j�ζ����-�'�(8��h�7��ӥ��c��Tή�Se�7���E���j���G���w�5�a|���`� *��&[���Wb�J��v��.���&�o���K^`����r)p0{�GdhK��r�����4�	Yh���3��.���{����6��O�S]hG�Q�v,�\����k����$YG�	$&�S�4؅a���u,�+���W{�4,�M�,�P���Z��D騱{�x�z!�[b��)�T��h����J�fb�'ʉ}�����L���80Xl��w\P,�:�@��dCqU{���(	�R���`�Ej}>zƵ1+���!P(G�Q@���"R�&^���#������.��P:�y��ef�NX*~`�b��&z��:,�v��Ҿ��&S�i�
����>qԵ��8�H�z��>�B24&����ˆ�]f��K�=
p��c��Q���,���Sߥ<N»�`�'�q�2��$��x,����ͼ�y�u!$g���F��J�piv�Q�y{��� kph�e���}O�k3\G�L���,��%D=݂|#-O�M�D�-�{QS m(��zy���\�!C������0*�WChm:͏���m��%�E�㝚��5T�Y溃��>�l{��;W�,�H;y/�TO��T�e?��&�jb5��$��u(<�=����)Sϟ���[�sC�)���������JK���N�ζ���SV6'e�9���+-�u[�F���h�-<T%�"���:h	���b�q�)���'XA�������
FVGFʇMpc��ˉ.���卸�(�c���:�im�:��1�;���h[xڡ)e[�ݷr�v���0�^��i�fc�ރ�g�A%����n����-�4X$=�f�$�tG{z�7�ƥ_�E~X��C�ʗY��L��5<&���v�s@ǌ�~�QS��ט�ӭԺ�ė�*��%:��!����?(�!P�p��=3)m�X>((�'1�Mz����o%�BquT��9��g��LC�?�X;Eu�d��O���Sa��F	���6�<��xZ>6E{z栌���p"�����P���V�t�<�e�O��}������5�=D�ǝ6��#������O���G�R ��5᭛��dk����\��Y`����S�>˶ǰ��vA&^�ȡ3;d� U�-M����!�Y�O2�}���� ���*�L�ch��߅���Wa�n+7��D"