XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>e����:�߬l�������b&(�D�c�wၒ�˦o񭾾�v�|�'�&gRf�ظ����#t�����K��<M�����Nz������H���r��&�(3�c�t�/��2��������k�$���X��M�|�W��`�Щ�JMPl�����/߿���Bl�	�v
����Fnk�s�Zz�� +�T���p���P*Ii�N_�&5�%����1���@�JnKr�����9=a�zP�OVr|1��#h�X�p-|����l-,$��;F��1�L,�����{EH<W�|��w³lϨ�Z��%��Z@P�n�mZ6���눉t���t��j���a�Ʀ���#^�p�uNī�D��G���Nπ�jRP�C�-)����n��i�>���B��KE�7cj�{x�����bCN��vգ5'�%gc�=[1K�� k���h*	�.Ț��dD�y���65w،"���8�"�y~�4j2�4�Ȩ���Ѿ��Q'-�$o�������/��O]5��(1W-%u�b�ò�qkC[��Y��@�����S�Ϳ�gTv�;nS>G/� c�y���|<��j[*��j	�\`<D�����(R<�+����"����u�>�Ʒ��F�g�?%�9i����ӯ�҈�=zz�����t��<����l����]M�͋e�d��b9\����3��5iꬬ�30z�`��Gx�g=�]��_]���xx��^MA��Y�0�-���,@W��?��ez3}]6�XlxVHYEB    fa00    2470�q��`��J6�O�+؜�M�q�
�T[+l
�FF����_;Z\l����b�����k����A�ߕK�ޚ�P��U�KN��/x9���x4�e���ē�j�F�ҙ��)x��7@[ub#����TA����dzͤ�lf�@�N������+@>���E�6>"���o���5�2HYZy]�H�dy�'�P/�|��M+�$ۍ9~N#���'���9l�X]m�y?�K�$�L��cV2O���yh�����|���y�b���[_]Z�>�b����R=t��w_���k'�b��˛�+��`>�lV�aAĩ\��[�AF����@k��sO������=�bH�%{9 �cv����F|�z�u5���:3d{���"�}�į��5| ~d��SG���g�e��t��lj���c �&?_ ��XP�]�2I�\�P�� ��S`TB��ɯ�*�]-|d�Y[h�v�a�;����p�^��2	F�� ��֟-Y��/��r�l��tO���p�2��\H��/k4��厑P��bu?�|�&�Ն7�k���@U4�>-UԹ����2jc%'�� ,�kk<�����OMg�\X�6��֩(��y��Q?�	�eW����|m�M;��spEc�o+&�<��3W馇덭��}�o�DB9�n���^9����o��	���m$����hX������9�G��{��vQ���ƻk"�{�U�/�%��?htĄ��=G�w!���ʾ��P���b���u�@0�m��/a�0z����/1~z���j���;7��ZP(2�u�f�O
G	ɇ����$�0�ړ>:u��Pf�Ԉ���1�3]-T�zG�"^YfF'�B8-q��.�i��7N�!e�j�Q��%r6��>���YtV����<�
�i3�s"ID��e葫`�}��)���@۪0�@ ����T�ݹ(x��F�@;�W[��@��N#��z�a|�T�zZ�~I��ݗ�C6
�(|�Y�A������]��w��WM����<9Yl�9����cOjٝN���Z�����Û�[�f�߸�#v[ط�aP���ր�b��R�˭|d����i�֞]�X_��VSv��H���ji��ZU?-�'����6��������Z[��z(No��{·�bAu+u�3ī�����\Y�Wǒ�'ݨUq��fSޅ��@ʻ��òH]�����pW�Z���j��mB1N}�!-A�I1�ȣo�O\��6c�m�I����v�C�>c[��f���"�l׿e�9oI��0YR>Z�@�l(&U��}$#����~A/��*��R������.�9Oԍ=bDƿ�+����Tp�)Z�8��H�$� ���ָ�Y$F϶n[�%�z1���E�$"�r
`z�c�#� Jg��c�|���̨|ϱ��N������j�$����P2/߉��o���4"��+`ݙ�����C��)G9�I䪻b�'�o��R�@9��yeg�@ԈkO�#w&Oc����-Hh�����aZ5i()���;�&��uYEfnDX[�SV��f�V\���4�/D��Ez���Q�)9�66�0�B��������C����_��Ь��<�%_FDjb��<��+�\�e����S� ���T/`ta���_nE+P$+�G��A��o�����A\�%o��"�fB?ܛ�S~�S�ndd,:z8�~g�V�ʘ��p�lQxk@���
)|j�-���*<T�1E��`�E�)$&�`p��a�^�"s5F"��'i�����
M���W[������5��}�:��Q�-���G�r����8���ۑS�m����Q^?�A�?� 1��d&l��f��x�((#w� O����pm4�V�:��d�r�Mm��8E|��]�l*���T¤\�V8� �v�5$/���aa�Q��(�BE��v;I�;�{/�FC����\���м���ӽ���Q/�JH�]֞�V!�w �� �>In0"`/�s8�%p@�gR22T�t��!���j���Ì��b��m"�w�r���?��spX�-�?h$xj���G�̾cD�_
����@D�('�U[h�C&�щj��}y�Q���Ů ��֡�ɂGď�ߖ�*��Ǎ_���F��N⻎��o`�0L�>���tH��	7����j�40�k#�=��>*uY�+�k���P�FH�Ϲ0L�i���C�k�GB?:4X�[�I�rOi���5b/9�lAI�(s̜���HW&{�<�7��W3�� B���f��̇:U"��}dO�
8?���D;L�	�;���,~�g9SO-�ɫݾ�$���E��o�':��ei���(��kf��]�
�	Li�zO׋�����P���B1��G9�<>����&j�e3�4���C�;r�-��gp�
Ʈ��ޫ��20�j��#�s�+�y��H��r@��u+��ʚR�����D�39Ę�����	����N
*�UZ���;̎��OV:p�����O��:�AF�*�#t�����X{7���9��:�T�+���:�Q�j��"I*��S)/=�V�wʜ�=�a�����.��9�t�e���T(�&"��iXr�!F<>�����P�uV6���35�e|78��@�ׅ3�Z�죩����0@b!��XC��ބ'U0ȕ&t8�1\�G����f���?�e?{4�oV��QLݧS&swF�`Eֆ��e����)��*��iN�t���-6�FS �R$|�B�D��]�<��U�6P�yޭ�;t�g����X^�~�?���&؁���_}�U��ˤ��x������D�(��A��m��Y��%1�,n_�E���%f���(�����uI�K�)`�@X9��t"PTI*�j������c���!�8ɗ�y�W��׬����O���	�l��<v&����b��T�ϖ��/n��h'��Y+�c������%���➫�F�$� F�ˊU���h�lo-��'�����uΣ�0�� ���X���}~a6j��2n��!�g��B+\���T�',�?N����7Ɂgg4�6�:Nl�;�W>a��.G*~���I�P!�J�uܷ��6�>��p&�� �|!��mJO��W��O�:�$�&��*ZsE�3�d��F�g�7��HdD�g������F�u�.���@&3��Т�V����/͆�gbƛ̂U��;d�Ƶ�yL"z]��W#o)�=Ԡ� �aΠk����.S�,��!���&)wf���:F��w��G��Q>Jz�d�;�q�	M`e5TV���s3H�P�����`���:��sS$�~�������GUT�.=-����^����D$�SD��IP��)3�d�G�9>�B�����OY"�c�J�Х�d��GV�?�!е&읛ahpc*�5K2Z��	.�Z�:AD��m����ҎH��_�t� �=�jZ�gxY1R�o��C���o�9�b�^�H�LR���է���)�h�xR��2^H�k��:_4�)	J`6�����^���:��.6l�r�XcP���e�i,s���zb	=V
���0���j[f"@�~��߭
"��J����V�kp��O�VrчKS?�/�v���D��t59Zq�'��3兜�)���F5ߒ/X�D�vT�:�^�]C��s�Q���aP���ˈ�_+1u7�)�놱$�M�� ��z����m�� ��eiӡ��F�����y�Ș�Zv�J8��2j���T�6h\�4��/λ���,�y/�����{d�hjm��Y�j8�E����V��ZoT�3}�-���4�'?sXG���a ׎�2Q�(�;��^L�-D�g���qvV�vv�Vb )����'��^]W��`8���^��y�Wx{�'��Bٺ�A�D:�/��Ni�Mzc�n;����?��{ٮQ�e��j�������/���?h?m{^Rd|�?� �giƏ��D�U>xgar��7ی�-D�\���nQE6�[�{����lV<�M.�>~%O����w��VÀ&?�d��|�+��oH�q؅gE�~���y�a�֪�a:}���H����ʂ��,���-�%#�u+���-�!�L�)³k�HBǑvE`L�<&B#E�L:ad�k����H���%�����W~�1b)$���2�#J��E5� 9~)��A�I'�aj���b����7ϒ�-�EW�i����E��P��Zt�H���֨�CB���e�W1]Ѣz�n*���
Q�g1���(��{1�S]�$4�ɺ9�A ߌ���&�g>,L�YbX�[�U3���I�h�e"���L�m�=�+Ż�k���R����@*'(��1}�v�Hbt�F��;��. 8i)x9l,��u��n�����"=PZ�G�fFx�rG��������ӇV�.�nκ���ƱȢ:Yv]����A�Gc����a�ɬd ����J>&A�xK������i�J���;?�_+�h���|(D� �,�!"%*OZ&��Vr��o�L�����|�(�V�ס���������xi�����W��[�n��\��L#�+9%o�)8���q��m5:/�<4�UD���1T_M��#Vı��2tw��QS`��U�d��
�G2P��c���F��.7�{�#�<�$���k�v1�*]��DՓ
���f�.���~_��`j��U|nl3��qڬp��e%س7�4ÞKP�Br��.��5@?�#� ��9p����d�g�bet{�Sȿh����ģ�L�I&�s1h�UFR[�n�[g�D9�-e��H� XWk��B���{E�s�o�I�����ˤ�ɻ!ܖ���mw�t-Zz�x!�L<�'��"�+�i��A�})ǣ�Q�J��0�����;�x��OKI�A[9�n��Mj����3�!q�I��Ά�KA\9چm�+�4��|�D�S�:E͎��H)�(��6�j�<a�BLj�x3�3�X%e���X��ZHN_��Ip�B�7��.&� G����I:����Y�LމC�6d?�1M�ʂ�\|M$�=��XDȂܖn3�;/%��d�l,2��PK��B��yB*_Fv|� ( �m}�W�T���@Lۮ�(p��9"�h���r����l�ES�d����Q��j����l��}?�{�Q��_Z�(�s0�8Lƹq�����X�W8����R�x�*����S�F��/�4�[u�%IC���X+��@𺏖_(A*yɜ�Q��AH\2 v^ӭ1�c�٘��r�)H��NXJ.�lZ�Q�����4Sɬ0�Alb6�S��F�=��8G=��B�k;�D��ی��bz�X!F̎�!I��,T����m+�Ɏb�y%����F��"�_�0V$��h���*�eD��L&9:��o
�3�N&D KOJvM�Q�c��p�S2�e����u����IIr�%�
e�b�4a��U�%N��i�R!�y|J���r4M�ў�'D���W&̶3�zX�R;�2�-�%�F�S��S�rRI��߁qӪZ$�ξA]��p��	���t3	��b���H���|J��^��]^��"W ����V�u^[�+r1p�NUH�u��:��Z\��sސ��.~b��)N�e�t>*¢��6̭��J)V%�)?������4�Sߗ",E��2Rɲ9q64.*����2_9C�2e��ٰI���'�snih��Dc�<F:��]nE�k`9�?��K����c�=<�w�`��-Џ��[jM�qq�q�\싘,�DoYz����P��m#�آ,�J+�"����Y��j�a�(_)�c���c#]KB(ߦ�o�����_�MR���G�����>�2���|_U�B�<�3p=�l|�����Qa�����<�����).*e��HZ䫭1+�7q�4mE�	\X�:�����Ŧ�� �qO<8Ǆj�c�B�a0���mO�����㫸3N�Uê�D3!9�&�%y3E�P�N�dT�Y������s���k��F���7���

�=¯ڰ���r�9��$!@�Q�]��e��B�ݳ�9��9�I����C���^�O����1�9���FTo��1'��Fp�a��ub3G���դH��{�AT�5H

�� ܭjY0�}��u����p���nYk���}�q�c\!a�W3��g*@'��\�@�X�Dj]U�b8}4��W|^����h����(jr 	��{v��DO�y{�������zڏ�[v�~�a�z}�Z���Wt�k�(��C$�(i�e6�q���Uo��H
�����/���-oX����@_�j,��!Q,�@R���߭2�%1��Q���_��w���������}d�יִޗ��"��a"?�S�:�OQc���	�ڄ�&�9L[J��,���]�10�\���@X�Ɵy�	o��(��� v�U+k��jΕ}��c ��	w�e�FN���3!�co�I�>
̹u�t߬��d-|�Xȵ;�þ��\٢05i@CL�n��+���L�x#'����NҰkC=`p�g�$H)�@f������4l�uE͇5�z�'���R������KkQ�뿟{B2$⇐0I���h*E�g�6n�V�9b��^ť�8]h�0�rE׏��C�����\|����̹w�N�0��o�m�ܖ��e�����kA^�fs���U����8��+��fd�l�f����,�6vV�}y�cЪq����L?���4�C�l9��
�_J_����^�@�1���dB��M�nb/��͎ �ҵZqu��9�*�z:h�lK��M��q=(�d^�$�g�麭��D��&�C+"Y�,�Z��.��D���4x	���G�(�-������FN�⯫�X	����=O( ��([{(w(����\a`�9�Qk��2#?��{ж�)e��N���&�����+;:�)���p(���u�e��9}<˃�PX�Q��� �e����A�6�¿Ky�]�*�6�`d���H�0�[2�Jc�2��'"v��!{ڗva(��*���+��{A����FoY�#A1����`�V�补�ëPE�{�������� �6c3m�
E!�3�� �������|��rM��~��k�@�9�%�cF�`[K��ϫp�u��bPJQ�1�1	ى_���Mk�#��U��RL�����d�n����W�M9��X]kȠ�,�3�F��~�%A� �>�
����.np��%�c�����9������h�-ӫ5�C��}�u�ӆ$y~*u�`Zߺ@�����0�々5���}^�����	\ �JW8�"~�t�N����	�����X(��Y�⟃[��U��Vm��W[�q��QQ�o�$_����!��HY��F�7�o��l�6'E��aȽ�݈E�D�\�!�
��	��N��X�I�5�F�4�]ѿ���$��i{��m��=?�ۊ��d�3�wTW�@��'�*��WC�����bļ=�H�f�ɍH�*$Se� �;�~rң�����('E��W0\7B:��d7�j�FL/�ݯ���K:���X���n��qx�%ӝ���	,}[��U,Ps�u2��<�/�y��`���6z
��e|R~�E?-Z�W�/-�M�Q��`�`�!�v6Tk��jѝ�{l� aZ=����JR�7��ш��8S�ܨ1p�����==Շ*��N����)2hQ��z�ηRܚ�GDS!��A.��)'����5�$9���.�3��@�@��oc+�������A�Im����Qx���-E_��&�ڶZ�L��7�(4�Թ:�),��S}]u�r�����(.T��a�'$ʡg.2�Z^w��~q,�:�?F�4����Տ��d5zJ9\�����T���DR�CKJ�o�&�]L]����C�hߢK��3��&�	X�jT�qXwF6�z���s�K���ңQ�<[�a(�R��X�Y.��ڠ��}�Em�sN2n��E��oۆ�>�m-3w�h{�����z
=�O)<�L��h��}b��OfL���v����UY&�!��\���c��U�Y[��2X�/�O�[���懊&�`އe`��'pw���9Wn������q�?�l�ɤK���� ��{�ެ�_��K���(�no��)&�;�Ή�*(��.l2�Э���vQ�r��?sd�m/���>�C��ȏu�P�w��Ƕ�?GZ��gL�uT3 S^;z_�3Vf�m"�l�h"�t����k~ci�Sm��w\�]���V��]&+�Ӷٲ���}f�
mbC9�߾�
h��O�ڢ3��E��oq���G�L���Ҝ��/ԥ
a�4ɠ5yǧ��Q��JJ"��u�b��R��YK�+[Q�Q�)�g�?�-5{�r��y$ҘM ���Be�h�Q����Ix��ϑ��f�*}��qE�ĜZme:�-��@�Y��nУ�'8c��<�9��RZ�W�c�1#1�·�uX�ob���A� H=q�ݛ��s�)^Jό��&��7�I��Q
��6eO��;Z���������"�|:_�˩��BD��:9{03L_P�$��H�w�^G���B�����̍�Y�s*,�Lt�:����Y��f�ؕTFbO�:lf��]�UOi�e&�;�?»�g��G�:,AR2oih9�k8̰0����I��7���=�h��g2O�UH��0��"E�h;i��>�I��guO'9/��5�������;Z�a�oMZ����m�5�fsmϝ�+��|U��|��<������i��ѴF�PVB��U����:'
���d3C�褵l&3Ǭplen"��+����rPjl驲m���ng�LI�q>�K��c7�� ��\���	g�	��#e�l.�æ��]E�oS���)$O��6|>���.0��i�a�H���!}��Ǫ�]���U�4>�?�]2)����D[XKc�3>��q��Z�������:'���u��c_+��x���SC���k_��U���-꒬��`�f�6�ȃ�r�
����5�?��LcH��P� \T�M	�|��F��O�*w)2v�����d�m>ܫ���������\�1�g?�l�f�JIX�Pu�-��p�C2����E�:�;�XlxVHYEB    fa00    1b30����Om�p�g_��G�Rxl�u�R'Q�榑nYJ�������8��yq'Ҷ}O��k�����4�8ʄp	�B�<�s�}��E?J��Z �����k�Qq~DW��fs�ILoU}#≚��hu8�IA�Bi����|!H�� d���r���y,^��`s�9�K<�"�H��L$�.q�W�ű��+��ѹ{9��a|�Mu�T]J�ڜ�0k̓^����i��L�W�Q9b
�l�t�����ڜ�0����B�s6?��wؒ�QJy ��퟿��V>�|�a�U������dڊ(L�iQ���w����e@<�5�Y�����S����#� �9,�B�y�l�cP�����0E2_��Hpj�0�� Ym������+aW��cQ(q�$��L���𛞂�&�׆�N+Zf�^��(��5RE���j0.�BwhYb&�
�Rz jX<s���v�褟!�ؠp�1(���8�y�ʚ7��B��C�(�Yd��`Q0(��6]]D��|��H�nn;�{�.���`9|���<$�]��q{�J�j��]�����/�I��OR�߈�ږg�c�<���*0+/��6��
�djL2�ݾ�|)R�/�.'"0�NI�>V�8��-h3�VLC���7[:���a���G{�O��}[�r2�e��ldf��ڳl��6/9�)2[F!�B�'H;M90K��1��ua�}�]�緷�m1���8�.�h)_B^��<�#P��W�A���U���b}�툔� ��A{����˜�M1P�H��v�l@�!�u�e��y/s9M�Y�^������Y�)��͜B�қ/o�)KY��jn`��CJ`޺B�.8Ҡ_�x8��ű L�ꅄ��t�F{u���ܻ�j�[�1���#s�?o���W@)XG"�.? �-�-�q0�Pr�?}g��Ƭ1|�|�g���m�sz[�/�b�T�cţNQ��dB�m�ŭ~�I�ڰ(�2]�"� �<��!�.���?�`�_4��E1����E^v|]��������A�2AA�:��w-����놹A�|H���ڎ��>��oN��C�� *�Q�xy/0�J�X�opV �����3�vR��_�史���.W�����]r�둀��72���"r�+Jc�]9/�ɉ`�����V�K/W@�B���a�Z��/�ǈ�L�촄��۫�CPwQ� �b�Lۂ�sY+����>Q�m�R����N��րi(~Ό���}�D�D8�U;R�$ D6Hboi�V	�.��<A�,�5;�[�%y��(��CNʵ�w�[\(��<�{�.����s��U`�<&βnRM����@��$�k���*�b��f�6ͲC�J$-�5�B��Kd�)
:k����BZ���dFۏyc���o�4��Ofs�|��o��=��Oh��V�A��\
��ڒ�jh�fV�������yEc{�	�e<u������KW�/wi)��׆�!j�� ���4�7e`�"	��p,\�j^�Q�����Ep;{1��+R�o�a��aPIv6ެ
_f����� �+���͊s0-�;�<K�O�-�Wb?�S����R5��Sǁ��%�)Z���	�*�	���~����vB�q��4�ޤ��穦�W�s��XZ�S��T�񸏕L	u���nj��_EB��YH�ա*��d�v����1���5�ti)�T�?%�����.��7R�K%���1�$Xp�p���bO�bsLM� ��M��������Z�(�ʺ�fL�/x��(�[҇�1�7t��D�����d��re��Z��l����o=�� ��DË���U�s/����%DP8��8�ł�xR]L�.'�|sc�X:��䔔}Ek'�_�����1M�B
9fASn��� {	��ZY+�'C����>xdW�:L�	rE�I�����M0����2�5����h߀y@:�t.�J*fߗ#q'���a��?�K��7y�#گ!�����(Q߿z�(\�ծ�LQ5y��$'�9��J=�T��ꆶ��ߛ�qS�)|\�ȶ�c��f�VP�Xkdyi~�S��W9؀�z�K_Q�r��)WR�p�=����mwTX��`+ 95�sX�!�\�������oCFY����N+Nh�:t�����I�P�_晱E�p��2@�0WU�B���҈Z���/9���P�+�� A*<��芽���>A�'tL����$�mp�'-�&���Š1�����!�,5R�����,z)�(.Ԙm��&o9�S0���˹���.ӆo��/m���Ӂ����0B�O(���ye�����d��S����/��6l�ꨔ;����H��@���>��:�����z9(�
�K��B���K"X[�iZ<�d��-�O/�1c̅%��H�m�<�����q�1�)!��g���������7�\��0й�jꉚ�p����Cߡ���M�B}��S+�%�c�|iL��(�b�=%y�V�lM;�����V-Z:��b�"�X[�ͨw�_ϋ?%�/��(o �w�'b�>L&{����.��� ���kuL�#��=����s�
��%��G���� "�X���pq\o^���4�
P�;�@�3J/}
�ٱ�ʆ��|��I��eXP�C�P�U����L��M~���]���өP%T�V,�5�������D���JC�YF�\�b�#U�Nߖ_�v�^��Q^��oф�lr���^!>�~��|B��+�r#d���s{?.UHf���p����혊�q�c�Ț���-����K�+J�^�L5hi���|��=����q�}b�S���� �/F��HD�)��&t%)�'�@'��n��/������9GO�H��uI�)w�5�EE�Y���5�B��	����BU3+_��j��?�N�ف�,���II�c�Eʳ�Y��v�{+�'o����ީŕ����������ד����E9�Ύe��\��;��,�4e#-�������9\u�ś�\�\l�W�n�`�$f's�ǽ��M|cM��kQ4w�w̭$%~��ej�S]e�OX�����1|Z�&��#�)����w��WX
9m����&�(���L��ǲf���;Y`��g{�bGp� f�g�u����P�[*����lv��)�zs��*SIt���G8���j�g�g &Mt��q�O���xPR�}���z|��=[�[�,P3��%uƵ��p_�>�3�ںg=`��s��V��A!�आv⚌#��^',��תX���;u��R���A���\���E�!�@���q*���Ҳ��$�O����ONY���=�Lom9賄z�{���e��\vA	�=@bC��ڧ_y�	���:Z˄�>��>�${_}���q�k�QW�Ta�tZ����a1N�R�J��"T#����0��]����ߚXh�ظq�^H��KAP�k�8���j�SvV H�LX��ʱ]�a��;�3�uݎO��jhd.ݖr�N�G(ʧZ�M��hJ}F��N(ro)����~�b�9O(0���k���l�"#����W7�0�Q�Gp�)ۋ+��H�XQ@Ѥ��GH�ad:�k�؄��u���+d��Q���@D�T���V]ͭ�!=M͎�	���v�b��L�(���*��u�j<e?�tm�jgA� 7�W���A��㈚�=7����m���< 3 �z��l�GI;��D�vP�c����Ɲq+nd��S]%�ljv�x�e2[��3+�t#�9`=$L�
��{�O�[@�B���sжI�p��oP�9���4�\d�\���GQ^���t��&9o���f�B�eICW�!|�p4R�ޮ�F����GKG���M��N��Wó�Quݡ��_�̵}��9O9���Y��]�a��S�p�u�E��mId�N�g�xT舒���qq�`viq���I�]l(�
"���<��o��<0j�RLcG�-�d��iB|̴T@�V��u�d}�ۀp���
h�"�ģ��|�]T�S�9$��^�.�f0�^��^S�3.~��4Z�В�'f��V���__<�1pC5�&�V67jl�tP�_���kEt�E]��L�S�)o�a�ܞ�A�]�&���Lau����;�A/��f�%�J�^�Q>)iޓ�x�-CI)�Fr�^ŻL����J͖uJE�f��vD�?��T�K�{�/�p����~�1U~k�x��g�,q��]ٝ�b�L<獍�(]�5Q�r��Y�VT�<0�E$���C�4c��+����]/���C��'���A0Ǘ� ���U�Ԙ$���m�l2B��9���c." a�n�/
e>j�D�Vke��컺�f�����4)�J��Q�{Jd�U	Ѓ�^	��٥�������9��m*"��[���П��ԓ\���b�t)~����O`P�~���_�o��=�Z���/�ߥ���e1:�u�ߨ���� ��@O��?�S7����T�Υؐ�}1�§�P|K#A��K��ԘrS!}�5]���"z[���1�sDJ2�Q����3n2�c����Tj���^y��)�,e@DL��&���@�L?d�7�>�v+�~���O=_:Xi����{>�9��XuL��梵U�xr�H���O��v�E��8ĥ��p�~���{�G��7�?n�ư��js���mt.��gPe��Ѹ�R�F1v��O\�Ȗo�8a�?��$T�+ ��96/�`�A�!��s�=�fV�X�Bw{X
R��&��y�}X9X���S��$�z ��~���Ґ1�|	�2��:E����4ͫ�z�	�%�+�~�V�nj�Gs�	��ߚ��N��j3���;ݏ��w�4���-!��w�k8�L>Jh�aq2"R,-�@�R�$�ih�,w�Ӏ�&d�P��r�T	���{�T�'�n��r�@e���94�K�_yy$>ژ�V1���)�Y�Ρ�?N��&�}9y�u�Tk��J��9h"y����{}�r���6;�m;��<��Ptf49��lcQ��+������M�"]xE��������.� ��+"��	���G���Wdi���!է��7,����
yֽ�.;\Y:^V��)!-yNM�>���w@�s�"��8OX�011L��<4#e�mߗ�ڦ�,m��?�;M����9�!�Ⱥ`���f�K�Y'�Dz���	��ֵ���H�U��<W%t�L�2"/Ɗ����EjfiS��K(�j��mO^�!�X�M��A�\����§�B�'Y�oP�&0�<R?ڿ���4�z���S�*O�{�2�E����@��=J�:��Y������#�
��hK�������>�#�_�ld��pu��&7��CK���:F�s�2���܃�ZE;о5_g@n��n��>�7/�h]Kj�4�J�C"C �˒�"q�.��+��ݢ���
{�F=�DɼG�(E�~6&	��8-�����
�רV��`˯�f>l��ZđW���+��ί��m�%�=���ԉ_ԡ�'�\F���$;�b�H1�}�^���5���x?�8]T�ݧջa�{Q���x�ȼ�>i#���T��)/V�Gw.��6��p(3-k��`�,�SZ�a�j�|W)�'o��~�يoI�L�x��2�'g�h��$!$WFa��^j��M�"�F����ɷ|���������n �{���q�F4�����e�߻���^��[h������?;>}~\�݁1�ϛ�@$W�L�BZ�f�YI=?��V�zd�rY�,���^�z&X~�0��+�nzmQ@��g�f��O�su��E.�Zo�rͼG��'�R? ��)��U���{��K��2�l�M��TN���2-��J.�Rd� ���M�6r{�����?-���o�9X߱���w�iw�� �����("\z�w̦�����Ź�N�n'_�"miZ�)HD��u@%��h�ʃW��յ&^�华I��i��=�z)i���U���=@��B�6v��i�y�o��J��N��.E1_�qq��@�7����=w���ٷd9��K�pC7�0.:��3�SԂ����B��H�<�` ���)�g��Y"�e�f���W��RB;��i��m�(�U�h�e't���ѧ�����9,�萴�0ҩ"�?���֗oOf��<P��-'dy��٥hO�泤�|�  pӠ_/�IN9��l���c��w:-z��^Ѡ�+�@��(�-��׵�K��Vڄ����[E�*p�[[�51�'��]�z����sU:��E�C�ONI�j�팸�@��
/�jU_1�h5U*}L#�lA[7~�4��-�ፍ%�W���P��8��I�R�&�Ѓ�<�HH14<� �t�j![�-�]r�<�||>��^����-6a\z���Ō�s.�S���¿�3eYR������r��y1�c�,EH�_H+�h���{�x͓��?E�_;}�p�kt�zD(D�q���@�����5�8W�����C?)T�Y���v|��*`�����V�o�e��JBg
r{�
�a��Cq+�	��@��a%�Ve�n�c]�f%֏'a�qp8f"�5ȧ������|��_5>����ݿ����ٍ�L���C�b�t�p�&�u�Iګ��\Fr��aa��Ѥ\������_� ����ɻ7r��<��J��C�3B�I*��̵�?�c�V�p��g�:���p�#��z�O2���>���}����i �R	K\h��NX�0)s~uR+N�Z�5X*���n�bda
9���*W���I�A���8��I��_��V�?5QD�a9�*�j�?M0>^��l�XlxVHYEB    fa00    19502��#�������*C���C LC�8�O�a,���~x#�Gt�)�MgAsT�d	@&,�V�Ob߮�+�	��X��0�����rk8�$e��/'�W�B?Z(u�d9 ����JO-&�S6L�f�ʹ�G�"ZE�}j�T滳n4��'�Y���� ��1�e��1b'�{��_�fdQ���*M�8�2� wym;^ i�?z�ژ�e�)�.%U�Y��5�㊟E��<�`�3O�.io�6�����R�C�B���u��VFlJ��������t$s���2{:8R��9䇷���T���O֋�8L��AR>�,t���s�"";�Is���C(�c��K�]��㱩C�S-���W�ƜǴ�b��{��B�o$̮�D@y���vf�����71GDK\[_qL�M�󉕁
�c�Fv-��o��U2�󩋥��w9Ĉ��P���p #��)d�X%b���k�w�YN,E�S��eIk��\�?VZ�/��#��"&��p���6��Xp��k_%� �y�2����Vk�d��l�@������^-�te>]�v�)qry:L��,^��.���������b�t�<��Q�s���#�����L�v�z"|dn���/�@���y�\�	�ݯՖ�6�a<u���)j�eQ��_l��Ԃr:�Q�
衜��0+�.c�NF���.�-��[���&����N�:�M$U�r���^���ze�S���	]�7�e�?��x��P��`�[�?�\����9���*��E qk�ٝRBU�Iѷ�P;��_#z���XV�y$��H#����)���ě��E�*/��3����#�W9^SۼO>�~�yy�[~���
���S��Yw%��P��+By��N-��g�T��Z������|�}�6�*�r��x���y�?*?ZR��G�c��E�]�-8� �ǿ.���*�"�&|�� H�Y1�)��eu"���6���d�B{c�ۇ�8D�U�V�����[�Y�M0t�!�R�ʤ(��64Ҵ_��γ�ǁ����p������.b-�v��:h��Ļ�j�;r��;%z$a�(�wI�����8֋M\�����^�
*WF�3*��ǌ�KE�K��ًZ��	� ц����iX��;
�����A�t�Fv�A�ۇ����'L���䕧b!��\�|Т��c@Ѓ�(�Z�&�.Q*��W�"U�����q'v�~ؘ8($6�	*?(���L$B� d�ym��62
��) 0�=���3��+�'k|h�����~���_4�KF� 固Q!��e�ݓ�wmϙ�a�Eǭ�m�N}�Σ��b���7���b�}�B��<�����M3ե�+#�E�]�uHJ����^����xě��8EOQo���0�
5�n5�|�u��hvNM����=e��V�A�滑�)�Vc�����#���U<O��� �����
�-��=��n�"	��n݂K2+��2�k��������ևQ|�ڬ;�n���c�50��UO%
���:�F�MH���>������ۉ����}I�{S8j�`FN	M��{�b)ω�r�Utv.��z�S�V5ʴ;9�{[-]	d�9X0h��5����3��m��++��Se��U���hV���6>�Eow��fɂ��fص�s�Q�*�`�]8�eP�E�	��y��rrq�4��@��{���q��M�TNV���.<m�v<����QW�U"���m�wsc>�{��oI͑.���ު�e�&4Z� �o޹�G:+��bc��ƅ"�FN��kfFL�z��cݸP)4|_cx����(�$�|R��$B]��؎�:�z������/`i�Rr�=��V��B�P�;��(5���wd���A�/��
X��{�)'�D���`U�Zr_�tR\�rV��7�����T�4��{��~ސ�DZ{�.����!��������'�/�,�y��ܡ���p���K��ۉ���VrR���Hy��V��y��Ie�DlS ׉��++*~J�_	���LAi�&��Ċt�����.8ю�Cg�I�6}����[ۢB�l�A.,M�;`�L�I�� ��рfh�<.[i,6��m�3�c��< ���(�1�ے}���A��ˡ�/ta�q�6��Ue�m#������k|a4d��!�!;��(:�d#e��fR�ǽ��R@�0����^�`����q�����\�{�Pg��#+{�t�qkwQ Q�^��4���5B:�F�y�G �tȀ.,�I!�3r�:F��7 =j�J�JVF��߬Mk�s�tL�AɋYG�����m�J,
i�L�LI[*"]���i���ˀ-�s)bJ��\�ǀ~,���7��
 w��	W����S�*A�WD�)���T�?1�� ��D�7��&e�FMm�ߥv)B^�� �nK�y��� �%Z���f���k;�oǫ=Ge�Ckm�������8ՙ[Ĺ"=��X=�N?���"��ą������>�m�頰�p5��z��>�S��%U�x�r)\�}��2��E�@���H䎒����S�&T�BE�TF`��NEz�+=���rB3<������n�'|�O�$P���'���x�gF ��7#r�B��Q̣yc+8㸍["ĠR~���MO�T	f�v��F!�:���<��M�@���LPe���u��1���7�L�U��*����.�8=�e )�úln�)O�)�*�й�oˇ��՛~ �@"+��V/F�B���i{ei1R��W'��?^>2��I��MTK��U �O��\U��;�(=[������#���i��AҖ�}���r*^63� OOY����L ���b�nb���L�!�����1ޠ�J�t����x��Yt�p�� �+)����������dS?�}��$l�U
w&�^�SE�'��f�U��Y�Y��.����(xŒ��2h�;��s�����OF�u�jq��"x�"VӘhDA�H4�5e'�����2�-�I��c�X�n�yA�F7��|HSئ>/� x���(�HM�$����: ���<w�+���+�XL�e�+�!���@� ��[�$\�/ӻ�J#�^��j����G�5�.�4���R�C�����D����b������x5�޾�d�cU�4� ���L^�l�>�/yG��;A��9�� ��AxT�tuT@\ݍ����a8�\��*l2f��;�5$�qn�\���,ƌGq�������E�$^`؆��2���)1~?��7)nߴ���+D�0��C(��fy���R��ǡH���&�JF�+k(z�]Ug�7N��-���xJ<[1>�'v].�(b^�KL)Ag��K:�oTHv��]ZF��S5Ʃ̓�,l0V�o�l�\[�yc�\����Y6��kYj�N����,K�z*�j��K����O<����<+�#���j$m��f����I�Ɨ�~/���c-�!寓��uP���zv頓�D1�F�C����U�v�Y�!�-���hֱe�mm��=&@g�p#x�i�������
_?���[֯��JY�g,pڸ)a��x`��6�������B?�-�{��$�D���y]�+�|z��[ @�V���c�����h*�?�B��uܗ�.1����#�=�9'�~-Z)4�ۍ�;묺EXM,.���r�LŖWU��>UT)>�^m�v�3b�����S
-�����7�A�A=�A4��p"j?vb�a���Tϱ��H�6���PQ��l+|�WS�����.�IM���X!^���|L�>�ZT��(U�v'-��k
PZ>:c�¦�)����xqTGʠm�����g�?`�\����>45��M��"ԯ�T�/q��5�n���c����"����V`a;J�*��&ʹ����	8=�M���|��5�6�QD<�&��ᥩK��=��wYQGg^ktC`�}*�yúa叁�#0[ ��f���շ��]m����o��F���duU��O����`���O���&�hL�ӽ��ڍ4 Z ̺���ה�Hn%��V�k�q��»,��.�î�b	W,�(2��8��l�O�7A��K]_�^揄6|�����oR�#"�%ʪC��A�n�W}2���Q�*����
���Qä(+	{�*�~��Y��#����a*$���G�D-���g�<�\���H���s�������o0Nv�nw��6",���3Vb%�ϛFp��L�
���7X�#����[N
�(�0��_к
z���9a�X���DA�e6ܘ	�PH��נ��]�b��m�К^��0���F$����0��̨B#az!s�|�jJ���	ӈ��'�'��x}��x��L�_^fq�����tt�a��7��·�pe��b?�c�P94��(M�o���*.��O=�DP��Zq�7h�u�㢪"����yU�e� ;ս���ʞ�9; �ᛈ��|@ꬻ��{�\�V��0�4��ޔ0��q�q[��nz�	�g�l��}�2�j�7#�(�J� �njUy�b���6���d�G[aޓO����~�j��*�Z�җ���s���=�l�e�f�ܔ�0E`��d-eO�G�>�ɏ���>��\S*. �ޏ�`|�,k��eM_�Y��0����DB�+`�#X8�	Nd��ҟ��k�2k)!:u�}�J�.�J�0;���#T�_�0&��yv��6���N���/;��o:i:��:7�5���N�����+����11�A�G�⫺��c�|/`�	���ns�jZ�k��
��Nkw�l��G��4=�u�!M@���[H�b �M�"�G�o�\�kD���^��K��Rv�jQ�L|İ�<��3_�S&�1�w��;����!�����݃�Y�h�q&�Bb��I~Kǡ@���/��ݞ� �C��l+�/lxw�2&��p(�a�:�	�P�V���V(� ���}�`;�L��Jt��dB�q$�N��Q �r�&R��UPLj
���\%H:�wP�Ma�-�bJq{,�u3��j�2&�^΍�)��*=�����4��)�#ֳ�4->�]��t�Gzt�#���@�p�0�kI�MA���Bz����o3��0�zQPij��O��c*1�����\͇�Bp��:�#�����Jy5�A�꾜M`�`�����à��z��τ��ke�n3�Q���+��[`b�
L�Mh\�%���s@Zw�-D�*�X-�S@�k�\I�#D99����9Uw)O�2˜v �Mܦ���sl	E���R��>�J��?~nL�aT��s,/�����q���7Y�I��7�2���uY_��H�G���f�Sd.��|S����1�T�Jw��q�w�C�(�"��N3������#�$��!`��S�WRn�_��+��w$�CT�WZ��L�`�pf#3�Խ�v�
�k9B�˷�i,�`/k#}�i�.V
�1� �;h�*I� u��tSz�;?!�>��ldy�b
M��p�a�<pxHT�_��c�F��E�E�8!f��$/_A$Һ!�$k���1���y+���%��{��)3
�z���Qb��g�84;!�����T��q3�%!�E��ƟG�˻ ��Ȥk4��}P̕�S�ϟa��1�β=�)RPN��0�m�<�i��4忏����GR�eKbT`8Y�]��å��B�p���HY6��E��YC�+8+�4+�{-֨�y?}��
l�hq>E^�t|�`���a��X��#�o�.����o����#fW���I��X�ph��oy����P`u��/��b�s��AŚ�N��ć�]��B�J���� rF�2����ِhތ�U��%�A_���� >��*ϸ�Mf�_�at\�ڪ+&�.�ʲ��^� �����1�&Z�]>��j�f��4xA P�(�@{ ]c�²n󀚈 tf�1�7�h��?9s-�����@D�<r(\Gm����� �T_o�Z��.�k�,�C��WL77�0������˄	�,�,�]"p덞oH7�v���lf�P��0D@i�ՍV�8/�Tշ������z�Ӂp��a/�f�/���`��p^q�6Y8�ND����0���+�3�����ѓ�o6?D\;��i^�t�����%8Ǉ"�H$y¬b�-V�g������`CR|�����_�b�/�T����d(���u٤*�$w�gm���7V r`�!Ե }�TP�
FuqWG�����y���W��(괗W��mw0�1�{UZ���dM�E�	(l"��$2����ZYX�q��p�svB�n7�(Ks�M�ԍ1A���J (���GXlxVHYEB    4f27     d40e�'�0a��@�������(������
M�LuZ���h�j+p�=W������+��W�_�UA������2̌��V����WAU���O}��N�q�ȶ���'����Y�ʚ������.J_�+��xa�_���[������I��Ps�+�A�):i:����d�.��)ּ?tT���'��q%�!����C$�S��M���s�w<�99�PNm{�c۩�:�1�-[�8x�AL�3�+��P2�V^I u�Z���QL8�K��{~�5׳E�*@i�J�ӟ��o%�i#�~H-d\�����O�"�ݻ��j�)��{�\��gf����dak[9��?�-S땎*h�t�$�{�,�s�E#���v ���j47;`w��a*��|/B"͡3)rF&�ͦ�������-u�R�1���� ��K0@x~.�VJ���o�[�����5iOի���ˀ>���.�ĀDE����`�B�L��>j���K�H��m�rcF���I�	(��5#�8�@�9Wv���Ka6����K\3� b� ���H��SW;�WCwX93�H�?e�͏%5�Ej��%v\��D ����/����|��ʡ�e5kg�<����$A_��I�P j=���^�$=�6�Mi���\XK�i�"�`Ћu��$�_��`1�ř�b���9o��y��~f�Z<kw��s�i��k1��h���a��a7ҫ�s ��ԂL�� SÐ�Ц+[���WӠ��q�2���A���'��w/[~��!Q7߭�Ⱥ�N�M��@D9�{�ڴ�\۲-S��$�v>2��b�r�4Y� �z�wA���̤�h�h�t��3u��mH��=t�eT(}S�<����?+~lDEzJ[$�wEdx����ђ�����팛>
*o��Ե���m�Uڹk�E��O������7>71Ma��;�� I"�@׀A4p�}�JsR�Z}5$w"��먃?XIK���e�b��h�#����l�֧ V�eJT?�����仕�kwlT�d b�Y���OC��#.�%��2X*8�R%n�}���~*�AYd�7����k��p���&�8_�_�!ƾ�Й���\B7�=D0�lz�8lCy�O���"|�c�7��ۧ0��q/�q�)�-�?ȯAA}Xɍ'-?l�#)����	L���Mi��O�ɍF���l�y�U{�z���ɉ�Ϯ�kݛ��
�Y�ꦣ��6ȉń�t�.;B�����q����7@]3���A�'�BbdKT�+��Ĩo��l�c#t ��8<��%h
M���^R�#�(�Z��@%_�+ ����j�5��H��DD��o#��{��7ۧyN,�k�
[V�<V��[�y�"AX��P�$+����%p[.[�X���Zm�4v�ba䶷��/6��2�H�(�!N�v�J���y�F�x!�أ0e�*qĚڠ��ix�(I�鲥%_o cǶ����ҿ<�q�][�`4?孙�H��Jh���pńڴ�.�5濭6��oB��yb�.�)�ݳ4��bȿ�ܷ��H�:���@}g�<��*�߷x"8��⋹]՛�r�F��b�ٺ����8���R�*�I�|l"�m�\zߎ��g�Q�K��z 1ed}-T��f])�a~�C�	�4�{�|_��`�Gt:�5�]c�\K��>�\@��'�_^��N�%�9�ݰ�#�r�rAv`�A��}��8�/9ne� ��b� ��ݫ@����Wl����j���un
^f��-�{Xb>v�*o��.���i�pz}�[�4T)�ʬn�G W9�]�Ֆ��� ��y���h�e~`D\�V�}�&I��[��$�����^:}�<���{*S]B�xԐ]�`rj	{ֱ?��<?}FA�EU��C�x�}ٻkG�����o�h�*b���eE�V�r���A	0'Q/�C�<�w.m�hO�6��T>�r���Doft�/�'}ʣ���|�OS���pL�z��f)?�_+��w�W�;��C����ճ�W_�_��y>�ejm��*4�jM���D`k��8=��n�y��z$�IeRi�_��ݎ��	��	B���t�~M�$���ɘ�6w~�+�䴸��j�����!�'V�a���^��ٮ05�r �~��x�!-���F/j�P� q���<��A�6�]l�6!-$�%܃�&lM�2R�D���7�T��4��P1}+ˁ�> ����y&��'2�]ç�o7�$�'����;#�L�z�3	=AFR�ZC�/o����w��\v�-�ʂ1=e�����&���Z-Y�!�h(�6!j��K���i-�����r�cu�/u�����1�q��r�ט��p�`xO�.��Ӫ�vߛ#��0�Q�%_�+Cn���n�-�s�<��������5��Z�b�8$��L$�����Ɂj7��*���;]��r�1k�w�~�����kuW*ڒpH�kJ�@'�G�v�6A�rf��|B�j��*�1���DDm���0v8[�����х���1u��C�ӭB��f�myؓj�R�]ш���ʋ$�pfIۜL�Z#p�Q��A�+�&��ˈsH��u�#Be�P�U=z\���Ⱥ��͎݀���23xM(V�b}�H�l���&��&a���ΰ��xx�A_�Z��{V�V˸��	�J�!����ח�w-l�=��nsǵ�Մ�O���9x�t���[T"���2�
:��i��,x�pxF6�����;E10�ZHlA�FC������_��������!>x��f�QijƹT �W����5e�����W�����5��o�Bn���r΅j���\g;m$)���u��1��_gP�_*	CCD�uUDT�Goҽ��lU���`٨�bȅ5u�z V����M�#	��å��j�;Y󝧅�SL�IcN�����G-/�`hp�H�?���� \|P�hx�����)�D�����Hc:TB!u����I�����L)���d�+x2�r�S�^FX�B��(�������q�)����=���G����a���`�#0���3��Ҏ^>aQaL������,y��C���
V/��[��B�h��#�M�&èn
8[w�i8~��Ű �P����RD�%;ޏ���@�����e���"��#�]�6 �ᢤ�C�ѱfQ���౸&שQ��f��F'
�9d�e��ֶ� �O��|$xċ�=�5ԬZ)�:���s}���#�9^�gTޑ0��T�0�3w��m�(i���>Gv�/���ǩO�������P �#���W2�����?Y��ؼuM�TL� �⑼ס́�R"���qJ�P�~>�Hw6k-*�CՃ��P�(�