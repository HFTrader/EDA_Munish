XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�eo����zXۗK���ЋbvADmep�B=B
���3�h��6����k�E�m�������Z���>Ï�g1a8�~^C���kh9�L���31c����j0�<�̏�7�GB�-r�g��t�*W9�2�7��k`�:�%8�Df���Ӣ���]L�f�Xh�<��\���Eä́p�ZS9�]s��k����x�<�(�0���.$�]^��vV(,�6Bu&�F�ն���9��<$D��e�79������~�yv5��9�6�k���B/wZ
���L6E�����^���Ya��X�5�kC_�,P����!$���
����<^e1�%��aˏ���%���T��f!;L�P��!�-��|���|�:W`#$�R��$��^�ٿ���ηC+"�a�&��<�[�2Aj��u��X_,��ϝ�>�]�/*e��l$M���OȒ�)ȸ���z|.)&^CX�0�o���H�Y��`q��R�h��جΦ���{�%��A��9�en���NL/¿��7}p�)���rUC�	6��[�VNx�8���d���M���ë̲�⨔����^���Y� ��3�LǤ/���C���0��|�<��Q$�/��Hr�2�]U=��)}bpJ^�_|�GDQ���W�r[{�m#)z3W�y�� �ˢ]�oj��������#�V5��$0X߄|�c�ցð��R�:8��E� �S��ߤ�-ϯϙ�S���g�g��l�Nm�SK�	�{�XlxVHYEB    6346    1790��(7p��V�����~��<䛮������߂�Cn��-ȕG�oP	~-�헱�7���|�z'��[�����%��}v�.s�	��9��"��^VK���n1���L	�Ef_�ȩ�6L' ؀l��Q`�����J<�2�����^��GHA��&6G��ꨦ%�J�
8l6-E0����}O�3x�?�Z�A�/�:���و�`o�0%�۟ɒ��빔�\����%m�d�����gI��[��9��#����Y�s3ydXH��O=M/w���&Ԯ������`�=	nw\�+��q���<�P t��k���q�o���m��:�1!��d��R6�$巁r��'�i��-���v�(�,Y�X,% ���V�ν#l�����q��jW��Ž�$�}DGuUT� v�<�i+�XHY��K�q�I+Õ���FO�1h?�Dݓ/07f�.�$�
���达�����`9�ݰ�MK��M�zI��� �g�j6n'�o㨛Vw�%T�f(�$�P�\uN��1s�q!��+�F�&�m!l�u�s��e
���&^��$�� S-��Q\ּH�����o�}˼��PȘ`�����r@��7&���"h �Y��m��W�Q����'K���5%�و�]i�OF�_�U�Q��V��A;�)�^�eYw���L��.7�l�8ea���ݮ��bu	0|y�]$���+ܸ0��.�2{�D��%1�	9b�4Ձ�z���Wn��åfJ���]���� �����^iM��G����_�D������J��kHX-�ѳu��b��I>�)g��*�dLF��BBV����=�[<��CP~U/��� ꢚ�+#�6���b
�;yyW�i�*����� �Q#�c߁ͣV��E\��Z;�|i��p�t՝G$F�Pӹ��f0��]j*g����}w)<�U��T��8� & B����ޚ�7"%P�춊s�n*qw���Nj�R1�������Ғ�o�e��X�٩7���Dn$���'�jx�35�E�~�>yߤ#���v�j�r.�q@���� +�"e�9�:Fd8�Mr�*0ëv��AzZ�
�h�ϖ�f��ˈ�kj� ��w[ր�g��6�7��g�ɼ[y�W�e�F0HQ�}���d�h��m�S1������T��z�d8@t�I��ۀ�M�:�V������)3�e/��lS�V�E̋�AYQ���T(�u(�p�(�\�{���)|qmN�h��U
*��f��l!׽~�!�E����.�����W�.z�L�����=����X�\.�xT'�ūFj�{����HT��D�T��u�+�-~0~!�$�( f�w�;�UTH��w^Q�9�N�;zi�6�ު]�����.&4w`wz������,�EQ	�|oڶ[@^��h�#;��E��%-����lM��j�Yo�{�#�Z�:�
�|V�܃�Ԓ�(��`qw͑�o~��8ּ./X�L�]$���A�
��Ie���8	�9̒�m_|��Y�h�$E�P���&��7Ed�Vf@�dT��k�>��d�q���sk�#R�r���_l�&�����ڃ���*�y��� 
e�B��F;J��+W�	��|V(W�vb�/, %����ۑ��:�Z���C�X7W�#|z���Pz1A��{+d΀r��흓n��d�#��Ԅ�o���:Ջ̃�u<���.]�c7O��I�>��L�6@���5W+�s��+Է*\K%q_�5$�:Z���*-�Y�ꄠ)4ꨡǮ�K'���J�&��T�4���@1�
eg5󩖕V����ւ�
�wrq��Ow}�R@1a;[�A�e
n.Y}쥿!��>��ta�[��TC��U󐘐����H� ^K�Ϝ�w# ��E4��w�S� ]꼑y�k����Q;���r;s*����\'xu`��Y�a ���Z�B�ڧU�_t:4�����R��U8� �^@����y��ADK�:�C+�pf��=J����ے�$��ī8.�O�4:j�P�譃��$9��1�>5�9��o�N����t�!��xa��ABs�_�<��|R��Z��.NJ���2���`��!�q���I�Nt�$������j�����G0��v�c5�u*Ux�
sЧ�w"q�)O��<8�B�z��F*_��1�
��������޸�L���2�_u�~��"�S���1X��U��|�Z�lY&��p�S�M�b�wK��ur���ר�%��i�c��,��Kt�Cv�ݑ��4Ws��.��ǭ�L��#��%��5�;��8��>k����?*^�({�������ϒ�(�����%�����Ϸ�",���m�(E��c����C�W��uO�N\8�=�QX�j��=#���G.�W�BV�L�'~�#�Pt��j�y*.��������%iլ���o*g� ��s���o��P͏sӜ��g�7 K��7&�D_ue�p�ÿ��_�|�e�p�.�:7�\���.�NZFF��]a|,��=Լf!��`�M��䆁E�<�� �,o���[c�*0���tiB��״�M(Fz�j;nQ�9s�Ŵ��Ѽ����x���~0}��:zE��,~?KI"@*��{���Pk!��pŘv�y5z挒�鲒�Sۥ/}��@�6� i�����=�T3�u��RI�qFʹ͉frv�_�+Y�h��N���fa��  e9`]�Wa&	�l�[5WS{.�h�!�fHc�s�(�Z�y���a	7��7��lI6@4dr�x�OuQ���<�Hn���#voʅ����M�+�3��x�gzzk �R�G�{������K���	�����Ң�X.K��k	�oF8�\i�v�|"��
�."Ү���KO ͂=�%w��X�<��m�ϝ(��M�5S��2È�aJ"�r�/���͎���/��}?���90:���!�5��{#�n'�i8e;���a��7H�K|�	��Ƭ�O7I�#�R��H��
��I��q�27�T�6�Ŋ�:�U-8�!��D�-A�<��ϔئۇgd9=�m@��eo����xs��M�L�m�nR༽�wȉ�V;� {�ҒR(��m�X�d���Rs�s��+���%gx��yixp%��?B����\w�[4����J���S��	�[V(�_*�koQa���*�e��K��hʔCek=�J�РfSA�8�|�3��I��QŔ�K�5�u����5�^D�u�KU�_κ�;�<�]���i��=9{� �h{j3�-ǡo�ӣ�xo7���:]1ș�G���L�����E�	;�h����
{^����^��nė�f�� [cN|FE�2\C&⑗�Fb��Y�������c�t
��D�&����E��s�T��D���Qpv�VlZv5b��R�L6���{�Z�쵚�.�A�����W�T�_���b<�BiQ#R�MŴ��<SXS���L$�ٍ8Ǡ`ܟ�OD0զ(��O��a�C1BZ����������t¾�`iZ�D7��<5QxNϝ(S;4��� (Aք<p��ŏ9A�m��#/�M͸���Q�v�Ñ�F �"g
(O�-}_f ��,��֘D�sf���u7C��=8�3Hr�SP��Mx�߾���CanҶ�Ƙ΃/ ��l0CB��I�R���M �t&�'�@h�	V����.Aiܹ*�"�?i�ǹ7�.Ĭۆ�+�Ēj�6n�􄩿�;JփFQ�Q�?B�w� h���RAWRj@�g̅�#6�j*Q���\dJ�pDX�\?\] pԔ��]��XMtv�A	�h�������ҁ=q�N3~gHB-j�B4"���r�qPs�g�#�3	t Ƅ70�NIA;O�lZ4O
�u1a�������NP�@������
��*.s�y���8< L;��+�՝��c�EW1.��IZ�BQ��8/�G��F��lC��=ݬ�;�c4`��	�&�������II�0��9ð����l�9v���"�'���OP4�s�>�+J��&QC��4#2��Ne4�Ҵ��@~[�2�l��* ��T$�ъc��U��dUr�1�$ݷ'm�iO��?Y�4��ԪF��<W)��ڪ���i���3舅(�v�ZJ�ƪ�Fc̥K���,���-/��~�vRJ�f�����i�� &��l}��l����q��T��ha�A��Qs79Sߥ�J����8�7�� ���m0N����]!����M(�PN�N�8Vf����9rɐýg�pG�p��gF�j̉��� ss*��f�I3>�����hϧ����MܚikFʦ��6���{9�(��j�Ԅ�a������bݩ?pnP������6?2�rͩ�],��y��U�,|J\��Dɰ�,j�613�< �T�9,ث�y���^�(�L���R���@P؈�+��Y\���¨G	�Z�s���V�R� 4/����{`�O�$�H�a�"h�LL�]?��p�ȅ����dq);\��n��8���kȕ���I�HxQ����u,�
-}�X���~N�AF�ܫ����R���*�X\������ �D��9F����	u����h��V���z�l���c�03mq�G�RN鵈*��\�PkH����'TWS+��B��;a��a�b;���z
�W��s�o�谘'�6C<�s֓�SNߎ���o,�@P�:�j���$�?0*˪b�B�שּ�i'�㳲����WE�igg���͵l��Gr2wlء[����[�.W�PL˟@���HL����c��ټ�ҵL���öy5�oX�{�-R+����*�Ʊ�?q��I�wX_8��X��` �����*E�a(��j"��S����9�Hg��'�.ґ�ϒ����9��L ��4l*���j��s��q�2�����Wѕ���4�x�R�K�w���=���LxY��F��叿����)L/�C�̒�ٽ?�]�\��5��v��1nv�\�U*���^�B�A���$ DļiH��hHw*b=ĳ�$��t��ٌ>�@�Am[����VYF9�1��1��;9A�������AZ�7|�#B�!�
�?	�p|�+�=�b�m���xb�0�$	a*T{��)v�D ^�y$li�Eo�Q08��+��5�*������K>�l��2P}dr���!�{Ū���hfM�}�d%�'so��Pp)@��P��&�����<�F��XÊpP�m��Q�wh,0DZ]�)���$��{³�{����:o4x�����k���$��a���H�sԴ��#�G�YM-��i��A��4*��I<7�@4K͡2h3�W�W�Y��ςx:?/ȫ�Q���D�5�T�]AQ�_����"@��C��f����YIH�x�h�u�/�_Bg�+�W�K��Zv������e ��4�)֮:�m��n�W�ḑ�Ü��R�����K�'f&FX9��x�.k9%E�Q[������ҿ��s����?��'mi�^��[\<@�t#�/�=����ݯ���?֊�oe6_��/8��]�����$�����L\0m���#��*�c2]/�29����/n�Y< �o�2NU�G�j2�_y�C�ʭ�1����f�,)�%%��e� ��!١IE@� 8DL�a���n[�Uǌ���
2���2~���� xq��Ö/``�Cf�Y�	��sx-B@�x��$���b��i�ŲK3��b�PJc��f�w��NN�<M�>��c>4�iF��ۏsTu?�����1Y+ChƂ$�lVy�ǌZ��Co��R a�Y��ƭ��Q������p��/أr[4(��g1��Z�x_�ĐWabVx��m��Ωk�+���B�Р��	m���v�(Pa�C:۰�z��X�Ӱ�Fj��