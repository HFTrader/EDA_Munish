XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~A���v�4�q�Y�*Z[�1/����C���ہߙ����ӫ��K��~fy��&q��v�ܳ��^��>�{X �--��T4RvE���a�T����CB)���P&�;vL=-r/��~��ͱ�?�Qh$Ή�v���F�"��X�Z�f��5�FX�"wlޭ�LŎ���ҝ�%"�!�b/«��k�.,Xg����c>���"
��\U)��j��Ki`1I��f���k�!��C@[5��I8�@^��y,�����]
�#���I\{���ь�}x���8̆>��_5ycohs�9����xW0$�g8�����������|�ܻSx*�"~h����{d��:�^M�;�Yt�A�m� �A��(�� ��C�т�7�R�xJT���'����b�U�zr)�&T��5�!ѱּ���׹��m﫜���0�w#w����s�3�T:&m��ƚx�����]�@�������f1���k ���d����+��Ӣ:~2o[?���]p'%Ab�K!��=�z��S�<��~��e.f��F��l#	O2b�����'�8��IR�ˠ34;m2�(~2��#��i����"1<EL'��VT�����􍆲�J�oi�������LT~R�ys�8US�]u~fK-��3�G1?��Շ�fH��Y2��r��ASy��w���-�q�;��^٥�y������:�;�5݃;_ܨɞe�D��CY�#?�\�5�ףR�-~�XlxVHYEB    761e    1770S�9�ٰ߇����ԩ�zBv���A^�j�L�� "4R7=* g�������r���ʱ���1%G�|n� �i�V�/<�j��!�a��;��)?�)�",zQTy,u� ��#J0�z,����lJ��"�̷�H�$%V4��
v3J����d���)�;�W���DL���Ҡ�7��</�I|9>�z��Q���E-D�'����D��z�i=�w[i�cw�7�N$��Vw�������M:��+{�6s.��{bXoQ�/�5�WN�GZ}O
��U��[�tBB�[���9�N.��^�%����M�z�	}�@X��ct<��k��q� �v�ka	Z�%�I��:�E��>}��_,�%�N8�Ft9C���𺈣�rO��[�KX
�U���lZQ��%���g���C2_ӈ-���<�[&w|�rm�6�)W-��qc�r�v<9t�A�����W�
{����̐� ��$�_�U{�Ѷ+!h��SU�Kla#�m�x�?������iq1�� �C�Δ�ц����љ6|}R
�ar��k
Ϸ\T��_��)v-�1�#ܻ���G�y��W�16����*�������l��S�����#=���|ֵ&}X���nO��3�}��X��-k�G}&1��ׅ���@�g�-0�Ѿ���D��J�<^���Qux�e��:�&FVFB]�����ܦ��kճ�w@hF�ƜC�z��刓��K�u��A��:�7	�Ca��=�OS��3��lH�TwڔDMJ��FC� �-vpƢ)�<��^R%���.h���* ���u�Rv����S��c��*��%�P�ܝ+�q*��Ք�S��},�P��={Ē��сո���2HN�^M��������&�+�}S>9��Ez��<Y����x2}b@܈5��Y����������Q;l�q�>:�Y[��;ރ|�g���P��5�p��T�*B�D�ʃVG<
r=>r{ f�,�G`ޘ|X���_^3�K)�b`޵(4�x��ɦ�҅���Q�ςz�M����������h���������[�"�ͨnP�Hw@�}brMy�:������b��=،?��U.��mF�;Γ�{���k���p=�
}I��k�H��"|��~���v��_����L�=�@x|�O����c���Y����H l�N��.���xdu:�%����n�w��0f�'���F|�tY�t��vd�^?	١�U�>#�W	v�h�����^:H� V�"��|my���L�	��x�D�I�nLSJ�#4���5Vhu�*���b
Z���_VN�48�m��JPa �<�ũ�R��Ҥnu�.�I8_�L.�";�k��BRa� ��d�ռ+�-Yg<E��I���9ݒ:��ί��a�)l?��- ��G���_��l��H�3�h�v-�GB�*�$[,��$��Qp�K�����f�ۍ{7�/�2�[z9g~YO�)M�Mݱ��~6���� �+OŰ:��.�	Lt�g?8�L˫b@�	她c�>#�*?��#�.
�G���H��Y]N�*!Nf��=�}+J�=����3n��GZ�7�_~\��eI����I0Ӳ�;�\�h4���!U�U���HΘo	.A�
��c����6'"�g�\������YefV��k�Dd�R�!�g���/tu,!4�y��雕�Y�l��������v�s�%X=���/?��8G�@�х8� �ʍ0@;�gi���N@��" �z<\YI��|���k	>\�.j��"�T�����h��f7Z =��;ȧ��Y��j���G��$M���jA�%X��6<���:����8\�U)bBq��Z�a%B�`�����"��JMd6{�0j)�7�����ͰJ�ExT|�񗶻Π8��1�E��r���V�pG�O��D��#�s����/��RCIKc���{�˹b����(�?��l�S�����F҅g�����3���{�Ǳ��?�B����{��a~�g���S�P���c(Ä��0���ݮΧM��tX�����՗�en��#ɼ��$��s@�;���l�|�	�~7D�p����C���)l�����1�t��?�J���$Y
�(ςw����$Q�;�ح�Y���04��j����hC���N�©KRcۧe�DA?�B�]X|�޼�Y#����)Q�X��rN���J䌳7�X�k� \�=;�O�����j�˰��0���q�����O��SXŮT�7/�`S7G�#�m{`�����.���O�U�E�)i��^��@nb�}�@�BWB�Hq�C�INV(�C�g�#VEF��eN3����r�W���!\�&�܋*��֮^����Ip��j�#�m`7�����x���fẌ́��ok�o����L���9F�Ȁ�H6�Mh8�:��`��ŀ9�XnPɧ�-�R��73Z�2��	�aJ���V԰7o�Λ��"j��;��oi7�?X[~�3i�س�B](2�~Y �)A���q)0���)p��F��.q=�ұ� D[����n�H� �z?���n)u0_~ۨ�-T��s����ƅ��Q���xO��{τ�V���ݿV�%I�������Ҵq�|����h��y�ӑdB:�(�K�U�Frz�4.q=pt-��y�Xr�~��"��S���D�#)U!:75MI;*�^AER���S�t���f�hDa�b^�v�8B�'�HA��Ǖ�1	.�v�$h>$�����2�8|��ҹw�U.VVh��#�,����.aZ#�[w����wx֓mF8\\)��t�`�M/�й1#j�HW}�lI0��ԧ�èk\2�Wv�7lY��p&e��W,"�)6��s*vt���QS��U�a�`?�S+���T��hb%�j���nY�8 ��=s�q�[#T��'Ir�G�����|�QA%b��X%��Bv�V�(����MH�a��ٶ�y��� j�i�ԇ�5V��B1��㇛T�k��|�T-�X��A�a�g�CqQ�`����VQ�9�A�@�ۥB�=&��/�tޙ��7���az}E��\��5�g��ʡ�=�E �{馗n���AbN֢@�2)����N�XD�N?�������jo_��keX�$eFB���ŕ�6��
4�2����-~�m�Nl͘�Q���^��3�F�~up�����to��������<DY1��Ҩ�)��C�@�;d�&X`����B�
&��*�~\�3d��a�����8�*�%sq�=5����~U%�,���dC�s��JU>{|[�'�Ot���@l�RY�Ձ_�Hk�R�e�urkH����|:�A��5�u����ˠ�d/="Z��H��A}�0�L�x�]�����h��ra^E�-w7H5�F_b�Ӝ5�Z#!هN^P��{�Rʪ��x+4I����U����.�:�9���ΖZ2�SV?�L2��It�/�qAQl�)�������'���Ѕ�J�7cH��z��zqTN���B[����"[և�/&�9��[�fk�y�s2$CM����Ng|�֒6�Y-�Y��e��:����(L���H��f��	�j$��oH-�����r� Ƙ�:��A�b�8P<�m !��Y��`��M�B>�Vz3�P�|h�·�{�.ѱ�S&U�Z���F��łz,�4y��0:KN:1vD�hO�:۶��
Cui*q��x�Q[,��X�-w�{��H�o��	}p1�o�-ʊ-ѯ��1���{�!t,:���4�j�Tja��2��>n�Rb;�ÑX�W�߅y��T� ���((�@k����m\(z^��:;���"�3W���6c��!�l�9^s-�d#�z*��0��)'C��4f�g�M<������˕>��Bp�9�B����7�
���*kJ���5�p?\�R������}���ѭ{���#M�|�tD�ɹnz�#�1�oU?��)=��:�ŏv���3�OV�|"�%����l��+ʹ�we����R�tF��9����2��q�Α�{]�`��m=_؁0�)Qx^��xax��v�7���(���Fk�:��d���#b]�م�:V������7m�Q��I�I��y�^�s�?^�|Z�F#/�rW*	'%�f��BD�ۻ��� �����9�u9uQ��QU^���P>g¢<g/;��7p��"�$x�[X&�fu�°b��gť*��i w��r8�e9�U�|�P���vpkٴ�} b�p��������R _%_��6�O����|�n@Z,FTǙIΈ�2��S�9m+���yެ؄r�˺v=��>�5��X賹�����ޔ��ٌ������;/�#q4����!t���,�J�j��7ʘ5�q�
V�>-��lkBn����Dl���/�>61W����0��'V���¥Lj��0u����o^P�¾�<��mOP[��V�������?��H��'Q�L�Sg�^\���v��O�3�+R6g�(P��ڝҘ%�i������(��@[�^݋���SkQ�"s��ڴ�k������Um���������eu�K�� �!q����0����%�^4��5L�s����a/X����u�՝Yڼ�4�P��7��P8��U��`�*�G� �OoZ;��p�[�]?�Q�)Qg����L�,;�G�(8��&�hn�/݌bV��sq}f-
�#ɧV"�Å�H�1��:�K4<VeE��*^��	�
�hO�)�s
ǀ�d:�"����"����~&�n�U�}1 �GVN�q������']y��55�y���]�.�3��f�'߄+^M!��F����B��|�M��)�7��r���P+Y3 �e�����FM��t�`��1�!��V�k3�z�U4���t�vRA�	��Q�	.��L^^Oz��X�~9�N֮���l9�/�E�r�`&�����D��/.=Ku�#��������i�:lR����`�s	&�TAc��Ap=�ґȲ>����%7�;�e��s�r�
4�<��ڞ1;I����h����W�[;Ȏ2���eH�U<���N!��?����pY��C<�����¹��U���#����8��J*��ɀ(}�>��]�c���Ӝ��Fǋ*	����+ML��1E��#S�z1N�q{�7��:᤺��*�ZnF`۶bv Km&����V�����%�0��4�|%�M{�
��+��\�ʑ�W|����zS?�u�&�Ԙa)Qw���2QH����X���Bm>5�<����E6�r�zO���y����,:�o����;�	�Ƞ�י�!<-Jz��2U>�5���$��/'��b8��0r5yxh�.a��^R!{+��(c���ꡣ��2J"�h�1��q 'i�QwI����O�x�1��}�,ݡ!��X�����E�@�9�pk�C���2�Q.�Q�0�K�,ˣ"��Y{�=u.* �6c��ݓ�r�Z/Gh��&_8PyT�@�1� ������)U9;��}�<�0{�L�P��Yg�V����']���_��i૒|����~z�$�U�g�qi����{�C�&?pi�I��"Q����Rv�1���O��l9���s.{*����=�����eP��C��q4	��+�N�޳췒3\d|:-�j�[����+�?�zX�NF��՟1�Hk��}[�u4����7�8/cd޺�LF��sp������c��3t59�A�:.+�dQ�u���_�/ߋ^��J �p��o����!�����To�}*e-}òQ"���z��$>d����l�lB���9I݀{j�{R, �Fh>+5�n�Z@���__�l
�|�(