XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ԧ'9�N�t��v�9����K�9͒|�R�f�hz�bq�g�	�o��9��96OpA�#�f)��@��9��j���zT���h��r�unVk�l���.�uU��mI������>�L�S[����=���T��a:�6-<=;h��89Yо�wfr�y�H~6KD�1MV�yRy5�B������ť҅P�墂�c�L+��A`yi][�ڭ�4
��_2�*a~�ն�n��.d�ǹ��[>yvDBvdM�P2<�Ѫ�YP�$2{�7��GO��z��G= ]����|<������1l�c�$�q-�P-{��D<�o���m���:�r�zc��{���w��z1��[��բj�5@�(�^������$*t�]�;��4��O��sK+�=�@��.0�&�u��l�����h��9��|-�������&���z�PDuI��B>�{�ع��L�"������t���x�1���E�]��em���p���#ǡ<�~�w@�Z���j�����31qK38�~����{koE"�WƼe���$Vw�f��c��Q{8o[q��D�I�1�F��^���ߌ1�8>2 ���]�:�t�?��5' he��G$��h���Lf��r����ly��	�Q)�-���k��=��� �g�����i��*4K�y��1@Xb!U<�%\џ�fQ�J;��2��;fe�t>�r�Z����	& �φv�#b����!9=&$���pwhN��6�-T���;h
,ƞ�n��xYXlxVHYEB    fa00    28c02���O�vc�v0�oI`��fd���صA��"������CHӅ��^�� �X��Y^%� ��N������Յ�1Dzc�8�]Y��2���`m�+���/�D�ߒH� #�4;ӵIO}"�w��C�L�\�_UG�_�ӥ�܍,Μ㣶�{V����G�v�n��겕#mPY�<��B�n�%�X�1vع"U���s�`��ba�Ƒ̞-��w���n2U�t���-�Ot�ꍁ��+�*��y�Į��i�o�:�����ZGKn#�Z��?�	���qw��gZ��i{X�uf%�^�1�h�|B�f*�1����G��\[n0�dY�d��Q���'�ʹ�0�bOPlL��$�`8i+�v�������p�x69�n��ކ�A!��T�za}k+��������Y���p|��ŮQj�p�(��Vz��\o�Kc� E2�ŵ�̄�U6�d�ճ�5V|�N{���s��͛�I�ʽ�e4c֒H�3�0��K����)M�=�E|�&�{)�#�O�i�XJ���2[�=�ȿ�6u��X9�:q��v6J�;c(�6�I#0H�;����3J���	�:���V�`+�1�v�r����;`b^D����v2sw����+�ܥ�D�`"��C���?܎]�w5�O<ˎ���,4���|��
�ۧ�(��ֲWؘb[�}/V�U��w��^`N}sP�</�5�v��V�+Hx�pէ 2�j������^�9���|��l����f.��lO��1b��]2=�4I}|�(,?�A���R~U�=�"&�j�@��POk�FD
M��2���!�����ɂ��c�r�����:
��9����d���l��N�6Ч:�Bo)=rS��M��2��^���YN�8�4�7��-&d@2��l�p�
3�iXP�;�.$�F�����\�U�z>5`9�X?��x�7��A��I�`GFغ�w(�{R
`��A���e�!y����Lv2����nq��6&��<{�:3�������(�ǈ) .�4g��ɱ��O��M��e�k�e�4]��;�r���N�2����@�J�c����^6��T�ؽ�S!���.]�<H��Ō�Q;�:ӭ[��oCS�c�U�F�;��9�k�����mce6E�,�+�/�	f�y��t�%#9i����V�r� z��=�:}�e��cD�*v�cR�$t�kσ��ZS�$� �D+��C0N�yz��'��;����{o�_6Ry��1C�"i#FG�jvs��4�d�%\`?8�9�H�pN<R��c���U~C�ϴ&
�)�6L��fԨ�#pI��v�5ރ{��8��J����y��%|�L�A�Yw�Yp|�>��N��W�әP�&�kt��tP�
Kv�*�q�?�O�=�Z�Zܜ�[�>�����9���zl�V����=��Fw�(lJ�s��-�"�8�|G���:,
~s�Y���瞤��ڽ�J���&�޴v�/��@Lƕ�J��i�NE��6���/��0�@뽀�g��L z�79��*�l�I$j�+����7%����gƋ��������BR��*��H��.u��3����6�X<�J�rX!�Ũ����ϸ�,+d�`�,�y%t`BY�+�~F'CY�H�d8q��s��!�@�T�zl����ř��6��.��X97:�T3p4E���/q�=�ܤ'�`:�g���)�Qq�x���T�g}��}Zw!c�t5��������oM6@=k�2�k#0�;8��jxɕ��<�]�9�L��g��74��_q_��-[嘣�%�&ڜ�C��t��2ތmV�րL��ݞ���ĀF������@HY�r��4�.��}����g/y�K��)I�������u�غ�U�P������ӹ�.(�&{�B�S�ŏD/�1��e�&�=�w�I�4Sm�DW�q2"t�M�͹�� ޸y�Z�!�.�F;="��o�Q['5��,���=#�.yO*8@FP�0�؟	����-�x���^�i$������t��4'�!hm�nZ�:�s�g#F�S�qS��Z�B���w��Yk����k�H���-�΍��_P8n(��`E�s�S�?�G-k���W�~Ci�3+0��oW6��IpN;O݂v��&0M���J�	0�P�5%6��wq������J��F_��b^H��ܵ�-�(�v��h�cԔ��kIw��lk������8v:��������&��+�Vx�7�1ts�C�%���E��1艭(������D���Ѳ�w����38 K��f��]>�?�>c�~ཆ= �,�nCiO%�������o�*�����?3�i�)�<�Y�r�1��S<�Sݼ �v�Ts�8�yr�R1r�dm )��Ї-��@8yc ��l���p����/�Ũk�[ț0� lA!����Y;K�RLe���ntg� i���Kp�����zѡ��6VC�]gh�n��h5ս��hv+�.8��m������y����I"#%{#���ADwOQ��4�٥�WX-	Z�����N(�e �=�ox��c�1В ѥ�7ߟ�����:�Q�s�e(t�l[`'k�̈kێC%{���;���aFxq�/�EY�u�E[�j�,3���XY2\r��v"b�b��m�T�^���jo�����5~�E�}�����+������?�nҟU�CZ���,�ϟ��u����g��E��%IN")���v���"gc�$��Ry��v�=J�����/2���ŲWq�@�V�Of��� e��id�BҬ�A�v�-�z��i:7�;]��3m>���[�C��Ɓh�te'"&��,m+~x�^�8@��<*��^��e����d����C��"��]�Ai��B��J3�c.e=z�Y]���$�ޱ�DS~��<ey��ũ�ZO>/�C�3L�B�NQ!���lfe�y+=`��G�gx$��x۟�6mY�C�s���Ǌ���8v:Ld��Nɯ���x�ԥ�W3N�%��}Q2�P�Vm�@!Z7��&�X.U��*O[�}5�غ�`:P?:8]$h���z�n��s��l��B�����l��<*����Į���yuc\�ȗR|�?4��)��sJ\���eO/�T�� ��ހ0i�]�pM+KfB�Ԃ��mv<X�Ȣ���~�k4y���q?a,�؜�>�i�G
+�#���?��ӧ��p�����I1?��1��df%$��"%� ��lBr,�5X��~#�U]��1���$��Vj�8�j���܆�"�I�b��NչY6?w�.��n�Ĝ�k�i��&cQˆti)�nv�
ҶE� ������!�s����8�K�F.��.�Fi��5 ��AM�N��?$W]�e�?���o����w�|� .���]��rl��\Xn��gz��(�E�^�%t��u{߆�5j��2"~[���s�%%<f��'��#Y\SƇH�j]��Q�b�B���bx����Q=4�M�f釁�����c|9(��\��~�7=Ea	�J%��[��S��~g �#Ӗ@�ӛ��|���j��9��n,SM	/������B6��^I'���|#�R*:��+U�U�X�U:��Yq�AC�x���Wp�6�D�/j�5/~�2����e�tL+6Ԅ�G��Z�x`m6�o9s����{�Tv�0Uv7���"�v�}����A(�h�WB�ce����93����[ԩP[*[&SCw�8ц\��3��B�t�p�M_U"�U[��N0U�M�<�����p��rym�C�� ��K�U�@� n�Y��Y�&�m	5�0pm��"�����Qέ��wӾ�|'	�m`��>��t�a�.H�֘�x7�6BC��(%%����O�ǜ��c��sF0aݟ���}ӫ��]x�e�i$E����ܑ�t�VrpCK�Xȭ��	7�_)��bsQqP�[��,	X��p��TK��o_b�n*�%*����h���u��L�ゖ$��<%>�a���d���, �H�Hj�V�:N�C��I�l��*�����W������s�\<3mZaZ���k�ąа��O�2�IZ�ns�U��UM���Y߾m�f:%s�{��g�k��\����C�����o�'*v=;��%_��Mj�]�G�T|B4���!�ي�G[�%�V��u��r�5@�(�.���-\ڱ*llUo�U1�K�뾄�?;3ϙ � ���������H����2�<?��5���anPod����f���C��Zqf�)����7ŷe8��+�	���ADY�(�'0��鬇���y��o^�wH�������~O��R��Kd��R���$�z�J~Ē�«iT��o��3Ҧ�Ѳ
03�p*���7�$96_�.�T�)�{}�In9�(t �2����\��h���<l��G�u%�U;)|���ݩ������f:b1�����Q�j���Ұ��|���u���;XE�H1�@���O���J'>~��9�fUP	2��gUC]2	D��K1��N�-���.Mo�K�ѓ:�"kUL1��ec���ޕ���˿ ����d���⋔��D�bD,���Y�g��*0;N�+/]��]�V�6�Ѽ�,�XX���zK�?b�v�_b)�n޻*L�� M�8�m)=�%s��՝GD2S1u�AA��]8���w�%�*]�M��l�¹X�l�-Q�;,n$��u�.�����+�+p9�(�U�ȑPc�H��YQ���n�s�aq�|�E˳tn(s�φ�)@"҅��D�B��	/vO<�}�n%e�2��X�	������I{������[��C%fjt8Q	�Y�_*u�4u��6݋�E��%@��U�D�U7��h���A!��
�i�wӍ���"z�Z<RMw��$U�i�`��,y(��C]iʐ�Iar��W��!�>�;~k�m&Ӌz~+	t�I�wGˮ3[%��p�� E
�]��XQrh�f�����Ƚ�
�/2����O�t=��	0��T�HI,ѫ-��Ih�*'�!�ǄHa^�Y�OQ8d�F����^�	^��mΰT��ڐ(��8�&qps�,����A��,ۢ���٧�j����/}�nBm��i.�,`4;o�����=}zE���w�)��y���.5+��^�S�a �-�q�q�h�t�+v��Im�C�O��**�V���R�ժ����퍤�L/�����/�2W~JŖ^�a�Q�y`���bMX�6oю:L<���>=v����AP��ӹ�5�_�m�qЫ�$����I}�gH�%#Վ��y(�P�7�5�l\4����8�����^^C�F�N�Їr�J��*��1�0ON2����b��b�7<4�C�(��۪�ou��<k+e�z�uˤ��ՅI�a3n�6��$�����a����3aco���bhe��g%*���n�	������0�]�3��[�w	ߋ3�z>X1��	��L����tZ�:O��F�>���D�N-̊�MF�����cH��
���\��I�x�j'�.4y�L���k�ܔ��+|��_{�<�#T��oL���,�,�7�y�j>�2|��n�~L�mG�u,��3��ple��{K�R\z����b�����V���xX���JK���w4̧�s!æ1y`�F	y?��	���X�������������Q�0�5��$��<��A�a�I>�_s|�,�d�D%��g��k�B]���3Ab�e\�Ll���~M浃��j	��%���Ġ@�7�#5���&u�4d%J�h]W[��u�˥���	Fa⼒�s��}k`�	�{]X�<2�)�kR�&�,<�K������5�c��$iS���fH�d����J9b�t�Knr�9����A���ϔJq2�9�'�|�WG2��2��;R�ȗ��Ԥ���[6��l E�akʋ��#4��W�{C�v�>�u��Y+?���lX��ٕ��/a�d����A����J��yX(��ј�t�.W*���<���-I�qHRCu!�����p�GG�@5��m��|p]燼��-�Ycj$�-���$�6��)�����)��tV�,�4
��^���q8.�4Zn�س:ў�z�R*���ˌs�i�\�`�,p	#����|�4��|���c�0�<W�Jۄ-�fQVՑ��i�p���rYOP������WVdí�zu�=R��&##�-���Ф�B�is��� (�S��Rz�QJ���檞�:;X�;�%n���k����.�Fe;~�?�;r,��ǜd[�'���R"������j����T0j�>��O�m!�p����7`��	��T+���$�Y���sGB�M��\���������ρ�I�48#ͪ�S�v��"�!�c��ǟ�����3��u����1~t]9-(C]��]U�)�e�E/��yx��J�1:Y�b��W��~#i3|�|���!ʘ�U��q��[.Oշ�5g�i����-��H��Q��A�n��5C��J,�B}q4���,��8RP��n%��A��~'4�r]����~����d�xFF�丫�e��T�ߗ�;ĠظI�fZ�V3rh)�04$kt5ٙ���r�k�_���J�y� v��${��5T�����4��b]���s���[���	���̞x�j�ʒv�p���jVq:mh�Je�S�a��*� <J���3��~��-ĺ�v��/�(F<qż��TL��`gI��0��Z��X8����l��-�ˎ�O�>�k�C����`�u&��rV��s�K�-�i�����!Ԝ!�ǵ�C�[�nǦ����]d��¨���g�/"�����Dj_�F�{y`f����r~�u��KS��	�#
����ְ�vi�[y.=�����fa�9u7�&>�7�hu<��v#�0A�؎Z�|�\a�0G�O�.Ǉ@;Hyb�fD{�-2�b�A�Hu��c�]sF��[_�LM"M��C!.��)�i6�`�[y��T�HV��Z&�%��J��C~���r0>�"��|薒m�-l�5l���Baӵ�;��S��� z�V[��8c��XXo����!)_���f[2JL��{�O����N���}N��L}�+ߝT^�����D�;y��.�\�pTd��^W�u3�JB�x�J��6DpqUj���� 7|O�9}ވR��Cy���]W�<�i�a�ew�cX�Yh�j�_�|���?�N�m��`ͭ�v���a�/_��j2?���rų�-�t&PD���G9{i��y��b<�",�r���7��|0a�0�~+%>�֚���R᭖,"7==C�dQ�]-��G�)���n�I�V���bd~v�_ڒ��	���-8S���,���K�h�:(��]�2	��
�/���4��	D��� ��za�%��1]1��5��֥��5�?��"m�uM�uE��G�;�u���֎2ȷ�2���c~#��V�4���'D�h��ඉw';�W >
�oQb�qc�\7���QN�i��l,�����Q�J�fގ�,B�gI�kd��c�]�`z�p���U'�BsG��kA��`f�2���,`3�G$g�d7&����l*Vu���=���'W@ط�}ڱ��[�gU���m{�&x]p�7Jb4�tXR�q/�ۡx͸�u�Z�WJ�.��]4n_��d��C�@L�J����<�<L0;����-S�1�X��Hy�G-0�����'�\�]d�V{-�ɺ�4�)n�C�.VO�Ҿdq3m��ұ�cM�\h{�[��.������:��y���C�XN��[�N�Je��"��,��s~���J�n@2���9@2���	���i榪ۚ����pz�ױ�G%Sk�͌��)\I�n�u	՛���x�v����I�(����s�fP�?��(�:��p�Io���RC�"�z��c��!P)��b'�#
�#�эF��f�l�y[=����K
��ù���!�7i ���mԡ����Y�QKdT��M��s?m�デ+�фm�g5�Z����,��J{�)>�{k���<3K�($C��>f8��g��J�jxgiȪ�L��ꐆf#Z*�;&�iχ��z�zDPK�g 䂔IM�x�s壍���(,"�|@���5��L�Ջ焻�ʸs����'�������})7F��W����=�J�H�f�[�V4���cq#3���k9�F��(��QP�Й�1��H|��On]i�¬�MO줶P�IM��!��*�(ӧ��m��l����59�&-/�e�ĉ�a1���Y�pS/���*'�2��J�ۊ~���=^���-�����{t�c�Xp4ớ�������>N��)��U�i�A�=n�쨟I�����h���D͑?	�T|ٕHLt{]���t;�U�O U�3�И��]�
�����;�a��D~/�O���񗰮����&�z�C0h89vƻ^(əX��!f���a:��
9�s�|4����uUc�20��k�Vw�x���Y���.��@�x�!�ȏ��$�SS��y�}s�%�?�8B5��Е��o�/�����G'��ѳ��깭i�Z�hXz	6v��m����Xv;q�@�ؾ��ks]�ey4\?ߓ#�T�p���]F��<x+ъ��+O��!Q;���|V��A!D�eެ>�?��	�$��T�+�0"��qod���]"�Z��	ক��Hx�j���>?�H'��D�l��m�i:�4�x����EGn��;��n3�
6���vS�7`��	#��r��J0*������9󉭯ֲ�K_�:��k��5���Ҽ8?+ti���X7i����(9$>[�.�U��f�������i8?UB��8C�%�;5#��pz��x�u�7N���媉sƞ�,����D�Fw?vfԟfx���� =��M{���[�Q����z]�Tn�{cQ�����s	U�C�����я��)/��B]W*�O���2�5S-lNJ�,���X����vJ 5	���8�IZ=����a�HGTy�XU��L�4N�d��s��X����+i�Z��N0�|�Z��I,��*�EӵL`���:�Kfj=i��;�zdE���vȒWcw=|/RĦox
�Q�{UNv�L��&�f��O��n�ܛ �!�6��K��	I9|3�ş����r�ĉ���wwN~�j�W��:�*(N�
(s�EdZz% �2/� �O�Y�����EX>R�vI�K̭�V���V�_�K�n�!%���
� ������2n֍kR�_>i��ѣ<��r_�\��U��|q��cη�t`z�ǋ�i��E�&�0�zJ�@���EJW�4��CoH�ģ9T�`7k�������wXdH"5���,@�e8��ӣT��*������d����<dI
�>�L�AK:�/��*��=o�ٱl���]�O?(���@�*��tFxo�UDN�>�G�ð����2���BL+����%��6�J�y�{�Jϫ�w��<�ǜ�����`[Jػ^7A�e�ie����VMt#=i�c�XH���#���]'��r��oOer����靊�4���d�U���z���r�Z�������/.0eSb"Z���gD���:����ى�;�HA1�b�M��%~'�!ܛՆz���'������<z�����DF���f�,�����3?&�*/�ձWUI.�G���Tu�U��S#�\�j�'�������˅�m)HB��:Y�d��8�(ߜoEL�7�N�fT	�I�я��,Δ��ߕA�<�V٦�bB��GC��z�q��2��f��#�NaUi4�OԮ�� �S�uϸfT�>�t��2�BS���h�u�����;|��ˀ��(� ���M�"e�OŦP &�*粱pN����t~�:cg\�(]�Pk'��J8%s���j#/Y?�����m#��%p`iT+
�rKnT=3�CL}g��Q ̈́��(YȈ~�}_��'��G%��4��ˉl3��T�=���E�4������T֖��f�)�Ds��Ϊ�:Ӱ?R�v\�ǎ�[�k�gVvｃgL}WbMʞP��=��i����m��){7Z��}Z��o��&��iU�����CQG̎0��(���s�i*�8H#a(��I�I/A�q����c�Eb{娖�wGA��^1Mkp��2���G�+*�O��̯	�\�%-(�ʕ���D�l�M�u{B[A�XlxVHYEB     896     2809/l� �Z�.Fõ��5�qj����;��Qp7�/Ob��ihQ�M<���MW��E�)�D[��`�?.w���3w]F�z��m�3��A25�wBQ*
�Cyֳ�B�	O�|y����K�FZ�	���'��4���G"�&u��j�ZV�V"m	C��6��@�/��&3U�M�zI�d�T��!N|� {j|��8�qs��ɲ���j=��'H��Lp�"k3��N�o��	�9�R��<$��^#�ۘLG�c0n�z�c04P��A)��uM�d��O�,����tt�t�S'`!>�W �q>m�jU�{ύ�S
��e��6X���ɦI��
)��(�E�کc�DK���Z��-Ge3L��#D���&1jACiM}֟�TY���hwN�/=�X��B:���Ի	�O��i
�J4 �E��!ܝۈ."���y6|����
���V���^�3U�i��fC5(��
����l�I~�p��c�FPJT�@9G����~ t?}3�b.B���.l�h{���3?�E5�9����0j����:h=@ed���8�ξ�󗥋Ъ�eU�W�&\��r�ZN��bⰺ��r�R�Zh~f���N��d��Ğ���\�[�ӊ�r��t7�