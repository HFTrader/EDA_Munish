XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���sL�"&3}hM�6�����2�M�|=;_��4�Đ�^�ب8�ڠ����ާ��8��U$�J���P�TnC�6	ꪃ�=w�^�
�z(�YZ�� ��g���B)�o� Θ��Q��)�Y6C�?���X����\*�7��V���U佔0�� ��lNT1/������6JI�#+s��ҳܭ�O[�dCbcқmtɾlџ"۩"O���5;���PH�*�b�������]�Y�Dɐ���͉pQ7:��l7��#��*vY[.cN�Dt|J[�e ���D���ߠ�v����\��>V?���1��ZCx�p�s!�ɐ�r�N��7UZ�M�����G�f��pfK
Fm.���;�_�t������Ң�q���;�ñ����9��8	����lb�y�5/��wKï�\r�w��/_���-oWUg5z	W-����P�D�p��G��9m6�z�Y�2���9��h�Ұc�d4�}���e�ZA0H(W��?����ąW���e��S��U��F�]m���mNYK��P�f�鵟�6�q8�Ćl0ahd�?=�� a��H�;Xk� �����H���^L�g��_�4WC:]�.$�J�nL��!0EFe@,����۲*ݽ�%��4�Aߙ���u�4G��gX���6ȁ�-��$��1z�x���[�HŴ�<.�>ya= ҧj�gဋ���D�����i��0����[*���M***9��˩����V]Q�`0@N�XlxVHYEB    47e6    10b0����)Į2�btt�(m����
QW�h�GE[��Q3�iMc���V�^	���Y�=�t�=�D<$RW�.���מ�����eG&�7���|��?X_�xot����x�B#�r�y_p�S�`���>�6J��.剪�Jv�mCd	�5�RK�+�/F��YTG�~�h�^}��O�;zcc�]�?��Y��l���nB�%����(�b�D��۸���C�i�ɴ[�x���������(m"%���XZm�vGX����8��:�|����ĘO�#��]�鼦8"�_���5k3Іe���!H���:���� i�7tM���1�#M����������݀�]�.;O�\*��P�6,�4��fk��
/1�t�Ҝ,���c,���d���H������|��藉�k�쏫�H�s.>K$~B���R��Ԕ/E� o��⥼�t�b���l��_�jg�SJ�%��^c"��~�N�A�����( 6��7fRK��l������Yt��34Y����"��j���[���*|��\���k7s���M����� �+z��\^~.�⩊+��1��9���Qmd�B�B�F�LA
��d7y� ���9�r��`�R�	ޠ�4�(b����x��+�o��[�O	��-�!��\�N��	��<H��1i��w���V�L��f�${�І*��٠���{��}|�K��̹��*ː���/�8�����kx�k5�C�^�u?Ѻ�^�xĘ����i(?0��"�����w�V���Ʌ��<E�4=���)��rTiڟ�OR��R]�#�[�����bJ�Aqu���<2"k �K��Q���1�LN^�T7�0�=Af&09�>#zQj:��?$�=f��:��X�q� )�X1~�q����S���e/�%����O���8�l��}l�{����Z�����>�|���x!��_��p�4�|ɸj����k9Y���*�m�E�W�c�'�#H�����b�K��]�9�@�,L�!:�m���im�!�?y���F"*\���<bn��Z�-�B����Dre�_��F��f ��ϥ
��vx����}E���cxL��@
x��~=�����O�n5^H5 �!D����_t���7�Ii�=4��ټ�+F��)q�!�U�F�B��mw��!�3�ǤL+9�z,����y�-����î�j퇴<�8_�^ｫ�'����wM��JKk}Eg 	����|�q��N4�^|yK�����o�=�pXe��y�zo�E����������$�@>>��*#}B���g�'k�Q�L�kƾmp-������YDܤҰ~��\Ҍ�uq�yW�����!"j�<�Pg����2s�\�$��#�ƦA����q6�+�po�d�m凼��i��p�� h��t��x+O?�t�y��lg��:�Q�/���S�^#�֊{�[�������6G��g8�E�K��WuG���*�l�H���;T��!%�Q�l��؊BUTA�&�$����ipyV^m��ys�ǝL��ύ����Sh��͎[s�Χ�A<^߶�/�~ǻ����JOW�����E�;RU:?�m嚛����}��\�����!:��,jWt����Gr`(áZ\{�^b���WL�+��1�(��No��>|���<�
\�1l����I����f�����:�Tb�(��@ĩ˖�dձ����i�?N'a�M��!|fu�J�հ�Y�o�q�&*��I�k�O|�U��e�����6�ُ�\���9$4"K��]�?.�Z$F���� ��tz��h������ƞ\i���@���nN��LH?h�bW ZTߴ^ ?w�2e#:Bj��N٪�0��d!�LMꦌ*m-2�E������{�� <$*Q�D�?����l��
�H� !*�N��`r;Imq"c�.���.�@b�D�������$�쑸�����H��" r;��W�;O\���2�hu{�L� �f�k��8�Hh�Ê��Bw�O���pQ�.�;�!�:������Sd���E��$�ƌ��7>'���ﳗ�w�w�*]u��m���jӈ����۹E\�~^3��.G�oɆ-�-�#Ԅ=x�<2����#f������W�P��%zIL��"�عd���z�Y��o#Pu%�Z�)g�ø�p�bX�_�b���t�6�vc��*�$�q�a^/�󕑏2�1�`��F�In�/�a�2 �V�v��;+�n��s��R��ˤ�yUUF�����7�uZ�@��oԤ4k�!�9��f2�"����N���F���:�p)�R��;߫�?�;I{X�Ϡ"O�gx�b����f�^NKs>ɀ	TЛ�q���o�O���+%r$��%g�����g�8�L��t��V�H����q*��ݝI�;���X�۬�U5��2#7����j!Th� %�YM��� ^�S�38�n޿�)�}
�M����&E�o�R��*`҇sU_�K����h�%��l�<>-��ͮ#0�H&�(�*ѷ�{�ԛ�8"����+�����r�*'lDr,Y>rg}!A �Idc2���?
@*��� ���7	"y��p���}�c�{$	XI�
��t��	��t��f�2I�&,����A7�E�(��P�u�4*�:�Q]I����ȯ�I#�w�w���^:�U�� p�w� x����->���pZn��!�O���x-aWG��sZ/�ټ�����Gk�	bmg��<��!�LM`�4�+�_1"�x������]T�#4F�=�_-,݀��笧�n�|�K��a�Y��a9> �M�`X���@�� YY���о-�����5�*cd\�9�:���1L7����O�6��N�$
��T�?Y��4w���T 0�8Aj!�8*��1,&kFn������3R`����tbG�%��ٔO�{��{�}��Z�<q͢�o��aj"���{:H��v��H6-%�q'�s����-z��u�䗟�wn���| ����2S&S��"��02)���[r�x�𑄺�����F��y�ꟙ�@�+Gm�Wh{ 3C��f L�(>XB���x�I�����,�Ĉ�T�YC\ r��d��b#�.�[��<���^�nl|���5a�d��jo�?�Lӊ)���t��C��(y�rr�rx1�UH�j�����v��B|l�('������	����h���2ϵ7Ύ�#�	��pśX�i�[o7Ve~�Y�04�b1�ͺ�J���}(,�6LI	_���5�\�m��QiN�5>�
��da��z�e]T'c��o"m��{r�C�)�����j�m�c��p��@����ˁ�\_�W!��1���Ou	!�'v{��!C{�Sv���[����.�g�x�l����V�6[Z��>F�B%Ig�V���)?މkf[�B��t�P���i�@�NG��G��r��ܡ�
o8�`i>I�d=��:7�L.d���%�d�0JX�ũݬ��bw����5�ֈ5�YƄF[k�V`|��eP��pI�q�� ��w%uNF (�W�u)�Bh!z� �����ڿƬ��������BSQ~E4Gq��Bj:7Dd�E(H��Ŕ�G&�W�8ʆJ�����|�4y�%_���n���3���K�S��@>�����2��};�SbnFB�Wi������U�� ���`�&
�=�~Jm$� da��]�-�Q�{�.:�z����%�	?�G瓖>�O$G�t`���ڂ&����ejN:঒f�S��>׀�S����	o�9�-S	P�FX��s�jF�h����lTu3X^��܋*��e��i-����=t✋ˁ���{K)~�h�3Ut��J\GO�#jy\/em�ᢐb*,ܲ�PQ��TnЭI/��]���)�k�g��O�n���7�D��a�% v)����ȳ"��9�;�ɈЬ�{K�M0��MP�O6؂ce!g�]���v�3�II���_���������+�tc�R��!Á��eX�E.�dw̉i����/BS��)��1x�n�:��
R��Ԓ���Z�C���o�Y�W�D�͌���u������B�fE�0,��v��,!l�[E^Y��qvYh��lL���o"LX=~Ν~jB��}+��L��{��oZy���;���i�h��L�@&�;u
0x�>�-����8P���0=R!*�W�B/���t5��C)/G�����[Ǹ��