XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����"�����F�7���Җ���qX8���p S��h4�3P+z~��#'N#G�Ą������%>�6�ҡ�;�]�PH�v�C��tǡ?��ۑ��7wd
��C�����󜌏�>-��:q}�����3a�6�4�'�5'ݮiR���!q�Yp�WX����Ѷ#����21A��6s.�����tbS5�����!rbF�}�t�ϲ�,ӺY�z�%�"b��@���Q#uXX��g����k�UW�eȤV^gO��4Z��2�O,h�ֿ�(�c�4�N>+�C�U�s�L�g��RY����ܾF^C@ncw+���#st��o���J?��.^�~�܈rd�/qtx|��D.ר�$�R�[@�k�R�T2��"+k�����Ç��3����:`��j;T E����uÉ�y	��la)�Z��y-Y@��m5baNH���T��s3O^�W^�)(���25Nۨ��;�;B�q�-��.m�s�%we(�w���vO��v�Tdu0<�����a*��Fc�͖�v� ~��[����Of4Y�F�B�z� �SJ+%�?�_h���B_�KuM�-������K�*�A���n�ߏ�jr��Sz����jN�咼��/�4�4���u�J��#�f�,��<qo�w�(�����럇}�r��?/1֕���ee�?��Ґ����P����v�41�d����#����D~Bj�85�B��dY!5�Jb��{��O�>��N`ǫ���j"5���XlxVHYEB    1ce4     9e016e��';@�Vgm�UgK��h����2��Ȧ�e�#,��rV�u����?������EviK("
�Cn��HL�Hj�!HK���[�~�����g��I�62����e�7N̦A�CO�����bM\�d�L�Iڹ�uǣ$����j�V_���99���#?F|#�;�2~�����C��S�U�3�WC�W�e�~x�"J_ ���'�W���Ԓ�#�w�s������kԿ�ķ�ZvQ�8�0/��V��XN�"��R<1�f�gZ]x�x��1|��PpW�7s�rw$��G[;��Ӄd[Q�B��q���/�Ƿ��ba/j��A�yö����мn5����l��ങ�^��H���*T�+^�G}^%�p̘ޕ&��|���y$xR�,��
����`�b(�X>��iR�Y%��S>��3��D	�q�v"F:�LFc$����4��̟���aAo~&���Gw?�慉� ��ߟ���a�	$zTB�m/H�mu�fP%D-#X��Ж��"<�Xx�%f�&�e�
�
�QXǣ�0`�5guh%������Z[��A�E�w�pk�X;D���5�	x��Nm��1�a4�.�Xh��o*  ��k6)�/��j���;��=�lZ?�rdRXp��U|�P6Ja{����4uɚ�m/�_��!��B�=Q� �$�ϊ�a��i��̦�<s�p1�-�T�K߃��"���a��zt�x�:s�/P�A5�vB4�5�JКb>,�uE��(��x+�j�͢�}�	�]9����(��<�OƠ9����Ȕ�v���l[8*���J��-`���3-��2�җj:���d8/�C��1�8�&�*��w�2a�t��M;EG��;/�ކ��`�\����n]l�<>�������j�OvM+sЍ^�oh~�����B�'���9�� `���X(��U,f�!����8|�K�>,�-X�G3�rd�B�|TA��a�sI�+~Cw�f��f��XY��S@o�y<{{H��պyI�N��*I�Ģ���/�_.��@��m#�?0q]k8�z��ӑ����{ڦŏS�A�.�b�Q�9��7ֲ�o
ph�ͻJ�!CK@���n�#�+-�';�����Wa�{��>^x�	������~� ��p{��e����������O�`�6���B�İR��Q<~MĠ_C5��̓�s=����i�;>88t#/Cx合���jw�b-��k���ٷk�ZrR�S,,�]\��E�d���x�,�5>�-	�Z��TY�j�JK��D� `��?��1r�A��_ð��qf�Ɓg#6h��"%@�Ā�σ� [A�׶ߴt��	3�u�;��Z��?��g9]���P`:9��	ߗC�����}��Mԣj+B��U^�*u�Z1/��/�[k�)�)#M�)yӻ "ٽ���Cv}a;�xCM��(g��@�4]����Kpb9"TIzwr�ќ.ĊG��D픈���cb�/,�K�V��A{��������cI��I]������Y���R��}.y�����;��/X�M��@�.3D>�KN���I�nn�?U���=ޭ�+��9!c:\i����jhG"���,��23zv���Ayq�Ҫ�}C�W���UMǷ�a�|�1����]���|�.���m^�-�H��a�� �����v�b]b��R�%�@��!x6����g��y��n]�߬���Q�7��8����OPq�
_�������73c�X��D�]���e���E �w^��3��[L#
��~c�;8~�q:��˲^�����r��t�s����ֹ�ܗMP�����5�{���*�f�1� �@�}�wB�?҈�� �����
��/ c�J�4ڶd"O�zy�i{�����[n	%��[��廹G�yǑ~��2"E�o���a���
<9�??-�錡듶ʸ��鼻����[-u'ܳ���~nHN�i u7Yo��J��=Ȼ���/�>�<��l2N1z>~M�E��踉����F����W�"g�Y�1��tNKh���·���˩,'��.��8�� US��k��p( �h��m�l.�f�>oU��.^r�>+/Ykm?�)bs�7YA���
�lr�qnH��8X)0��珶�9]"(�o2R���yF�Z2 `p�i&8�zj���J����a�T�n�vϕ�v�p(��c����� ^e`	�X���N�y�c�Х��~B�2��S�B�u�{��a%�D���g��D@
��X$�+	D��N,W�`*�zok�T<�'���b����q'c���%ng�˫�!
�~V��w>��_X�9W%h��՝�l֏[�+�l�'7����ƫ�����beJz|�rw�p�mV`)"�U���}����;��w��:�qϨW6A�#�|R���8����a�i��$��å�I xk�7�{^�eE8���*�o��?��n2m�J5�D=t �*���e.�����