XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����c}ʋt=38�SQ[�M��a��=hZW�� ���UL��"�u�F�Ѥ���UޑM����e��Q�z$�1��xR���^�γ������H����8��	��٬	2����W~�v�,�Pi�\[���/ I�t�u y7Q�-5{�\�2޴�w��O:�����2r����<
Jgw`xG�A���4�K^��� A�<S� �L9����P;}-�����\�U��uF
g�����k��ߓԠC�#CVv��~u�K�4�H�c�~��#&=@�� ?��[�BM����A�X����rZ�)w�1u}v�f~�y,�M:`�<�1�,t
�mC� yq>�L��J�A	g�)�:D���� )�R��<O��[!�����R����V���/��v�񨜢�i;�� 6z���h�^B~0ȃS��,^}i����Xh��s�����1������֘ͻpߓ���ܰ�8E��ыHW����ߨ���ӷ��������4�xb.OZ�&2Ic9V(W��"BA�pm`Ʌ�Xu})���Φn`�c[���l�vGV����qI�h������o�~١���u��yf`�����x�\�K��P��(�y�r�L���2fJ�1��6�8�YR�8���"�Bo���{���*��R9���[�Q��?Cɫu[�.��2�O��s@��즇��į.r�yӂ\������M�h�X�0��p<��'�Uj����Y�o:�l�N�������"��XlxVHYEB    1847     900h�����Ր.�Vܝ?�"�X����>�,���WN@��-Å�л�+$5S��V�JA�7miec�gr~F����EpM_b;`ܗ��1ժv���0ٻ$&^����0P�@��v����̋�I��j�(��	&%��g	g�%篅EH�!���U	���&�����`��ğ�#�^��<�Ad�'/�Xo# T��A�t�7��� 1�\�~ҟ�L���Ϲ��=����`�{V��ƿMٝ���9k�E���L�P��֐TȚ�m�ʏޏr��BT�[�IKL��-2�Gc�d.sv�ނO|�Y�$a�@�����3�B��t;Clꦚ|8~46�y�_[��,�mЙ��c�r����E�����R����?Cя`��~����8��ZXUU��5B"L��,7*8�sN��/m��mb��?%�	EtJ�#(���[��-�o�F�N#�X\cc�٤�娵����u &Ʒ)R�,�s�J��!����X�.�������B��5�׶<���!M��$�))ķ.��{cY �� �,-iP���`Q6Kd��b�|/1ɠ���5C�#�poĂL���%����qy�K7?H~:�U=J�6�z�+k�0��0c�>1�/�]�_v/J����͛p�N��vy�	�R�$�O�"�f�jh~��v�_�g�W0��CVZҨ�C̜&��@_�{F��`�$?�A�E�=o�o�jX�;�'-�i6_�\>����ً���ӯ�7J��d������WG@����� 3�(�������t�	<#eR���!Ӣ�⸘�ۃ��T��i{+֩�S��q�5���_!s�_x���^�0V�
�UӅA�~�vE����EeW�#iQMR�{��4*��,�.U��*yg(�"�����Y�!�X��Ʒ�cAh�x���p�R;��9�vt*����I%2�|���4ǂ�y9�o;��M59$����O>xL�4���V'`t�S[a,oz�ߠ�ٗ�r����4��VU�Ԇ�wQ.���TG*���X���p�q&U#M�I�(`@%��*_�N�;'>;�y͝�*��s���fT���C^| �`�2r6�t���F.%o`wKw�þ���ɇ"�[S��z��M��>X�x�a)�&_�C�>���O���j��� ����Q�Ɯ
�*��=Ɇ��*10l'�@�I\Z�<;���9�tf� O"�j�s����_ƝZ��w4�cU��p�Ǹ
X���|x���z o/��畇Z��r{M(9Y%��+��I8Л�`��O)��|�h�:�j�Ҵ���U�W�F)(4�aRI<��p:+�<X{��,���O�N��т�X*`=�Ʌm�;G�@���\lӏ�5^c��	t�y1*l�����3b՛� u���[�b�:{y-ox��7�V�e�%]���g*�q������=G���
5�ex�^��x�������@b1ǧ��_��שc��ꦹ��Pz:&l�_c�,�[����YL:�5�P�R#��B�e�J���}���������cm���Hv�vݡ�HPņ�:e$C3Û�
=��|6z���׺'� �{ԎE�n&saЧ.��|������P��h��T0�Q��g�_A��V5�I@"+�+�N*&�
L��g(a�^�.Ȫ��k���p��|�λ*���#9�ؾ�ݳ�2�'�lq�x>T���Z�4H>�oJ�.Ԃ�:��ւ9����+\5�Y:n�4+�W`0��][�M�����,�E8X���ѳkIN��/�R�� [LU�yAz�|�����+���
����Y!D(\l�����8O������m�ޑ�8�_��K�Vt�|��H+]F�x7W����i��8�u�x �ZC�8��m@��A�u�/�sXBe�M?���oE��\)x���>�	o�~��}�	�����~C����hnS�ۃ�J۞�����up<~���S>M���sLL��������=��ᢇ�Eŝ.��ή��	.h,9��g߯���mY���f��^���Yt&�rS?�v��ݏ{H���-��n��W�DPWs�(������t�v:. ��R�uY��I@�lf��ۚ�=P3[�Y�bv��Ӆ*c�7��6���l[Cԟ"[�9bA-"��V�C6�.�5��E��|�A��p�{#;����\2S�;��a��B_s-:�� [dKC�Ӥ(��u{\��L*��V����kRI1u�d�?�X��Y.��x�,�r�_�4K�c������7���w#X��g�Ǉ;���