XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������B���K�w���%���s�Cqhg:%7Sjo��W��k�!��?�y��Ȓ��jNA�d�,�j����U�������`�P;�O7��U���+6ȏ�}PT��m�o`��@W.SY�vE@?;=R����ĸ �q���q��+��#׸��`�ოU����I^��Y��n_x�0��v��m��| ��gf�8!���;q�V2��h5U��y`�Q����P��q�U��B��E��jX�H̏���1ou,h�!�X�v⦆��9�R�=|�a�wg�ǡ�ݦŶ
잠��@[ײ���[C��@�?R��v\/���fY�L�BV&��&X�$��=n$w���[%g����5�t<���e�rfD"���p>���S�a�<��^w��#p� �y:'��,�G������|�ˑ}�F?�2,�q�-��z��`�IU���edlX��mZ.�S����$fr�VDC(�t��m��ܩ5}T����cK(n���y�<>R-N?�!�E:��Q��`�s벣G��=�:�&�3q��OYv�z�5�&��[gc׼>�<��v�h�y��2��S�s�9h�/��dQ�}�!GY���}��FG�t\=�F����9�u�v!�
��Mls�Pц��ا[������c�YA�[�7U��<r=Y h�q��c�=Oz���u��3�J��҇ʗҞ�8�3�Q�D*f�����iC/���r�Q)� <�Q�	B��;`��n��XlxVHYEB    fa00    2400�	��&.ȲM3����z�8>4�f�$�t����#��1\{�3>��r��o7�LG�+1d�Ixik"v,�;�`[�au���y��Y�/K�4����l���.'�P5Y���ӹ�rM�L�y ػ.��%�E�{�iP�fxG0��+�W-�晸oső�$��&���0���wb!ng���ұA���b�����ܳ
���_����9�N�)쫙�\�U��m��Qlu�	&������l�vY.�k�KJK��e���~5�~&���,�����޷E ��m,����P2Q����Dӄ�t����Lc��Eɶ�#]6���Y[?K�L�m4�h�%BSr*"7�n�q̕	^��,� 1i���V�s`���7����ؾ��䱋$�nJ���{#0��i�'�>��=�4/��L?#�t[:@z/B&|H	�V���0��r]5CΩ��'�	����j,��%Pl[�G)nǢY���M#�7�\Q�ِ(R����n��
$� J%ΩmZ�`� �~[��	�#�Z�/�m���v�t]����f���C����;��T�5�Z�4�p}A}!6�ǌ���cSn�N��k���	�ڐ�n��f�w��M�p�3��H�i���Q�������A�S�9q�a���$<)�Cw�x��j�}�]����'j;k���k�q��J�]8O�;�������M�_IV�M�k����V)U���	
X`L�����z�Z( �xrZ��ڡ:6rS�E�PN�s���Rl�n���N��L=�@?8�F�Xz�W�S��\~�|���C�7/б�k)���_I����Sϡ\\�^ў�"5,,%��q�gQl���>��LC��z/}҇��Agrz{�4�k.qgP�=�3��n#4����fg��c�f��Ȉ��ߘ��U�V'lI�-)��[n�@�܎jt!� �X,\M��lBuG'Ӕu�.�L��@��,�n�0�7|hXToV���
U�S���~�g0I��gw쨃���Qi+�F���Һ�"���b��|���-\�\+�ň�d�Mk������u��}���f��^�7�B-��kСv��*V.7`�A�&�rj���
u.�*&��N+�ey�\[W�~��Ӳq��V�R�%R�s�
�d'���OѮwޓ;���0M��l�r>5���^�Tyk43��%��Z�!�)�\	��l�s��9�So��_���]�3o:q����-,S�a�>��:���㋑�-o�Ѳ�1�X8��BpՎ���5bt�1�LMyMb*,� d���Mh�N���+T�Il���d濣�:�"J
Ԑ�L�v==�vm�6h
�^}X��Et,XU����#�g�_ �n�Â�2TD��f�/��Tf�~�8�ö�jyc�����j������0`����[��L�w]bG�z�X�
U8K��眯�q��<OO6��l�0��h����/�}IC|�j#�6�U�:����M`��5g�2�	=G[�$�F����B}� ����D�M�m kr�;���Da���N�c�e^k	O��=�3���A�MHͯ>,"�Jy���\vч^�4�;�A�f�{��n�|@���70���yJ�%�H6��
Kࣂv�i�I7�eRU�9B�^���?�GV �@���s�YCRw�`?Q�!	���<��WH��r�|؀��2����J�6u��ٟ��:M{��9cQ�d�$�W��l(�B�8�ȗ]��Xq"�a_���wZV�h�V��!L�p,�FJ�����3ӕ��Ӏ�'b_k��T��yfTLny�۸(;r����6�V�GX4:�P�k�uZ�8���t���o�5L0 o7�HDj&Zak1�;�cTq���	Q`Ha4�ڠE7����4��f���e�������U�Ѵb�����]i�j �:�!0d|z��Qw�r'���uA�Q8��^���%,�j�a^׺��޷՟B�ʃ�I��Ft��¾j1���PAD 2_�<R8�R10D�o�	4J���uMB�wX
&�E�5�qZ���{Q���x���_���d�5>)���ء62T/ڼb�_`��A��.h̺��a�����,�B[Ǣ��a���$�Cw�/� p�t��C	�Z���T���+I3�*���>Ȧ�»��0�y3i(iR,������QT�i�,��g��$M�J�O�.K�D�ȴ�(���[㉑E1��b}�F����g�ڰ��q�iB�]��-��Z��;諴$���J�]`���*��&#�V(�/=.e�*�50�uH�Bj������=G3������B�� ���z�V��C]b�fR	��p�d+�:��)��B!��5�h��Z~E���x��I��l4����ݜ�����ӏB�!sӝ�����%�N��b�2af���b؋�~���\m`��ӄ�i� Y���J�n	��Q��]�W���O�#��������ur9tF.�u���_���������5���	�-|���Dp45s*��3~��_����М��7s� c�\��CX���ا���nc���`�.���Ke!����!�~�K�|�� ��h�h}��lRz���gKB���eڶ���1�8�~�$�]��5aNN#����k��ث2�?d4r͍Bb�����9�"��7"���1˙�5�(Q�K6��"��S�e������+:�*[��6�?�}���#���8�	�+$]�% h�/�Y?q�\��t����^9�q��V_�jCj��Yr����2��o� ���/�\G��,���(�,��aP>��_>�UШ�i̍G� s&�X����"}�?�q�ևIq����|�� "^d�Cj@|�����fW��RR�2ݍ��c��*;E{o�Ts�2jUײ �Eƥ�����X�W������P�H����u�&��x���,�3-DjT�����jI��rE�g����\2�IzJ�(I���c�K�f(K�_hw�>Bef�'�h�����lE3t��r��r��'��,��2v~o �Ĕ,��B�?�d�}�x:;Z%�9+oq^��И*4&:�[-UC��q?m��M�a̠��6kR;N,�э�åέ8!->��]�{D#������w����^�SI�l �JR�)��3H(��Tɩ�&�]� 3�&U��#�f������YzDN\G���Ѝbul�D��#���%����+s\�|��L@�ٔ�{h�Ԁ1��R�i��=*�a-��0�_��ঞ�42�V�O-(Lt�K�''��jo����r�$�t�H�s��"J�E �K�/S�Lg0o��g�r�i��)\+��ueĈ|�.�2��F�i��]�)5�t+��1d�����/�G�����RZ!��nɗ'�M����ÑUW�s;[�u:P{*�]S�E��0lq�vR���qY:�x�����U���Κw�Vd`L���C	�b�ְ�5�+d����
��\�z2���[U>��Z�{��J����f��{^�BW9���-�A���Y�����O�����M�*m�&�[�bǸ��`���/q�K\S��,�3�N��oI=�������x�>pV)e�Lj8D��?��:��tx�:���;T6S����a����<ɵ��� ���st�a�A��Tߩ�큥+B�`�S�{Z�bp��6�Q�漵fW̸��!poX�Y�z�WE�:��ٷL:�0�0��H�>�U��;z�^�"u��O��U��u����|��d/3���N���8Cc�5�n$����L(+m^=㬡�e��.l�̻Q�oM:���ۺ}�w�:�O�%�4|ᛎS�)X��:jV��
w)e�J��|Cf��s8�H�bSf1/-X�΂����A�t�-�� �yc�#1A.�M\:GOHxwD���ݢI��5�:�e
(��!�����BZ�1o{Q�nv�Iߍvn�����G�oЃ@�_ �q.7E
I�|��Q��=U�x�?�4���'#%��	u�h�= ?�I��� �|��UTw�Ʒ�_z���Zz���.�2��[��qm�b��OƏ�Wú鉘~'o�ޝ]xZ��L�H�[}����+s#m����o�Ǹ���#�X��w��'��D�~!���i�4�A�K^�5+��\;��2�+dEw�JG�����d��[~W4�� &�� X���×U+w�Ry'����W.��Vy�sj��Y��W�4��^�9��$&*	�uɅ�ր��k����������d�m\��L�C�;�یaf��H�M���,���J��T��x �I�=�g��B�f�hD������f�5S��t��9�q����\�w�
�pW�	X���nD���F|�鎃&>�J�ƅ�6?�^5��������s�M��?$z�x�f���G�d�*7��p�f��އ�n˺D'��>�0<Ɓ�_�^Iq��^���x}N���#+S��CX�������g���hݒ�Ws�Zg8cx���|Q�0�b=��@��G�RBX��fڻ"Fb
��qrd>9��-pH�,cƜ�� �4���`�oم�C`s�,�<�,?�I�ȋ��>�G����zU�x����7���S��p���	���
���e5N��/��*��|��/i?�͂;�=��������a%�	�)0�|�$c;��ع��v�f|��Df ��+�!"	c�H@YJD� H?�g��';�Rm�+Y]���Sa���/RV�G�̰Z�ɶ�8K�5�e��F�]$
��08�K����FL\K{gwtҢ���Ȝ�)�ͤi�#](�'�rvwb�~Y� ��dN0Y!�_���k+,�rbÓT���+��
�m���k��Qp���I��;����Lz�:�.��jǹ���G�27�FZ����嶢+�(��e蛾W��g�a�,/Q��Z�_�-�/�n+}|Q5?�� �eU�h=�����|�ĉrJA�$��C(���	=ܾ��b�-yM�=�t��c�r��*z�ǳN��،��~���\I�ҳ�VQs��Y���/���>�����atk�]�Q n��9�fY��>*�N���q/d��;����(�ې�Pզ	�4���3e�ܽ������8��x#��%��M3������`����.Z��
7�;�k��`�Em�b��0�������/��~,ےm�����)RK�ips�g��-�ܑ��e��.K@��2<It!y��.�"v���m5l�_�o�����\0!�- KD�a��R�/��w���C�k8
IU�5�_�:꽃%�?�'M:(�}ap0���J8�$��t0�d�Ȅ ��قm&O�~L���7���Ȟ�S��^�r�������E ��{s�}�D�FA[�4��`6`Y�%�U�#�t^d�^u)�H��ʞ�P��_.}�3�j�c&ʷ�?L���a��*7��Pw���u�>�,A&KBF���sZ"x�	ϑ?�ǩ���I+SV�\�k�D�陸={�*Dn�R����l�\E,ņ�v��C���X�i�'{e�\Ì����ܘM���7۹�`�im��/�%"�c	����?l$t.�us�ހ���9O܆�Oj�̐��i^�G���th$���\>TP�QS�5;Z� �Nfr6�CeI��p:_���,u���[���8y�as�"�qUj�����[;�+�}�G]��V�V����5H'�O1�^�͟=�t�FG}煶�>�ݕK	f�i�[Ӗ��杇�0����P�`�H�n-_�"�U,�C���"An��#�7 ��+�KY���ڻ5����V�0QD���g��6V�\��jf%4d9F�I� �A �����8FS$�p���OG.�K���X��(+a�<����������~�������(���r�^h�S��E=Sp�i��P�ٶLI�ۢO�3,��vF"?q��:[G��n�k7=���H�E�=�&Y���L�r�b	��3��^�`��t(�̉��Fq�r�<E����g� �\�L�_;�J��7Q�8OM�i�7&�ᴨ����5C�����zb�6�������$�vs�(h� ��n>Os�,Fa�n^z���%���c�_�H�|Nض�TB*�ES�a	R����}v�-�v�"�D�F�g�[FL;z�*J$����6�*.����풐9��z!U��h�P�@�Vq`�g>DGG����-�ИɗU�(�������n���+/�[^*tݐb����Sl�(�R�g�s����ަ��5��m ��<V\N�'��� e3���)�K��&n��Ǵ����be���I���?3`G������Q�N��,�l=Ue��7l�R#%"X��48Wb��]�4\!��
]��53�jS�	 "_��krS,0�Z�'%/�@1GD�=O����Wd��;�A��rh&��S�8u��Op����`�^�^1�g�5v�a�N�0,��yPҧ�)�n�1�����R��������<�M&����b�,t/��!��1eB�(Kʐ���Z�+�<R[z>˘��@�
�����O��V��0q���VJ^����y U��ٸ��*ֺ���6k}!�C��m��4�q�9��\��:J=��q����{\��g	;e\�{��X��?���1�����#v�m-�X$4?�+���Ž�s})Q��S��HU\5�4r(�)��#�}9��}�����_D���W���} �[{� !;�=��� �m�Ŵ���s��B�7��G����	?'�J- �NY����7��8XP��1���-�Tm�n�z;��Y���fc��p���F"rj``��t�D���̖������]��(���Iϲ�@�&7�F�"��p�ƈh�(��� �RT�wB�ow��5� �_�`�z�?27�(��g�^��=ٺиf~b�P�W��&4��J�Z�hO��]�չ�Ψ���Nu�/7�/
��"l���PG`��~�?b�$��IP:@)�*�KNHS4z��R&+r?�O�-P�*��!9*]_�		�uQ��������-'5C� h� �ÇE9fGVG9�]#�� ���EƧw����D�P���|jf(�_p��=�G��(�f~��I�@���z��B7Fl^�O|�ڰ�pC-���dm���HO���WN��6qv|�Ql�dGk�l�-Ąu{ N  �Qjo{�!m�:8y;�s��t*0|�1ȗx�iH �y�k)�E��|�+襝���,�>�q�c0NȦFM+K�9��ŪRý�tc�=ѭq�
�8���k��L`��~�Y9^��j@�H qœ3��ۮ�����|�J�8�e�Nn��5�[�~��$��7�bn[��N��''�k��h��ڠ�G��Y�*- [��H�q.v"������_��8*�)�Q���o]�����Y%q��_֯H�h6䖰>����zb�}�z�����Y�i���L���D�b8XX��B�ڎp%+��O����i������9�J<�s��7Of��Е;�y����)����&��W�}���R����Q9bO��\⪧>��>�ۂB�3dh
Xo���ʂ{��E��͎�E���EL�0 �����8x��`��q�Cn"�Q)Wi�v�.�Ƚ�W�D��R:p'^��f��5�Fr�񋻝	��d�l�HvY��.
e�!WLq��<�N4u6R[Y�jJ�_�S]6�C��9d�F8�}������y�n0 _W���%%�˸j��x�E򠷘٠{��A��߽-��pYj�\\�x�tDG���.yB{�B�Xm#.z	%��Mnv�
�9�A*�)�V�|D����(說B߹A����%�x�WW��b/�6<�3�~7p3M�I��s�H����/�'X��_	�-�n���%����3�+�U��(���k�:�$�/��P{��@Ԇ�<'�����)��{�ʯ�����}x�?�a
�зl�qp�B��G�3[g�Q���N3�l)+�E=�H�2%Uc�%�ms]�w����r� ���2�d0���E`;�������Hle
�nq����xD�����Y��8�B���L�v�WI�b�hvU���[|&f���1���oqI�u��Q���%��K�CX=�/֪�,Ά�^�?&�SbM[�!T�����y㪟���a[�j'7��]k1�@�75U
)qZ����y��-�,�+������hA-e,�t��9�.
V����gV�I7�~B�N:�T΁>���T��~P�_|A���ķ���Y1����B�Ay��9%~�d�R(�f	���gm�� �r�~�1P��4�\���,Fe�� :�ڶ�s��<�t���B�%�yd,��� @{b�l�,.�b'V�;/�Z��(�0~dǼ-�y'���L��o�<Pb69EI_�(����2�bL� �N鄁�m��N�UiD&�0����C�%4Fg[���rf�]z�$��a����뗮��dQ�V�Դ0
�i'Y�\yjo�W�X`�KϜ�v|�v,9�d��N���7��5 &�_�oK�/��
��y�U��_���$���5^�
�V�y�wط	.�deХ�������{��mSACA�e��)���4����~w��佊*�8�����f����f	��8�.���NR%^B˪��[��ѐk�D.�L�'f�K����7"ef{�@�y���uK��M,}��}����my�%|0�C�`-��}3��9������^��T,�(����v�5�4(.�3������Fi"t��Ŵ��t �Fy���G6�j�2���a:�["�C�:�>F{�(�O����-�T��jσ��6Ҳ\����D(}��\6J���,��/'K��R�,(�a2{�tY׬Җ�]$�r[dΉ1ƣ�i�2�I�����(B����N��C��X(vh��A�@�𐰣l�Ѫ��z�V�ʸ�?2B�X�ZYu^�!L����������1��s���Z�#����J�$p��φ
D]E�@�ь�fDE=�1:��j�n�δ?��K�g�~��Mk��E�jhzz$��T��˿������XlxVHYEB    fa00    1d20������B�Z��B"ĬP{�����+�cü^,�l��k����4Xҝ��]��?�{���_QD�ٺ��������/��j넢�	"ny�Qj��_�ֲ����J�^��0�R�b] j����?7�� i7�P�ĸ�4?8���§k�\4�O�̴������[4q�62�G�hw%��|�"��V��u!<�����\��J���(�͛�✀����Q��9�r��&I[�5o��y0��(K����_�Ɓ���I��}��E/�G�1�uJn��?��}�o�]NU^�N��^ܰ#��΁C4m"�rm嚖��?H���n�?�<���l 5Y����&��;��S�r�����o,�W���F�}�4�L��^9;��gf�-�
ݴ�Rq�d�k�N@ �N޶�Ċ���yy�,w��{�1(i��C�� 3"�l|�4I��Qh��<rn/�L�K��;8;�T��j�{��D Vw�BX4�P*��Ge�1�6'3d���^�qK<�n
�oؙ>���;#�mO����?8-h�{�T����+���`&�LX9���K�)��G�z���Ӂ��ִ	�+�'`c�Y�jl�@;"�`x�Z��A�ϱw`�~�)�����*�H:������)�����ޛ,d���2��\����\�Zn��,fU�u��;��@�ͻFsd/�x�6�Q�r9�����2p1���<��%�2�Y�*�D�B��a@U9v/��ˡ6�R.�oqk���}�9$�//.�5!-\�7 �WѼI23h(�oC�b��������"���᪾�b�>��cZg��je�C�b��4ҪF3�{�R3��Ot)&%i)M9�� 
@&U�udq����1�A���s���`ak�$ȧ�ɦg�8
N=�D�bR�3�B¢d$w�a�f�r���)k8�
��x}�0�S�S'Y�@�)��ؽ�+��XFN<� ��!��m�V�`AK��C9�O(�P'�EN�5l+��A�t�~����`yjY��wV���>�9�;no.)3/:�����4�4����d �RB�g:��Ĝ�3?ʋ?Q��'})��qFǪq��0�z�����!�R���.&�Y�=�Z�m7�	������:t\�pP�εnyL�=�Cf7��\���\ꅜf��o�^�-����},zY�S���'s2r�L���P�F����_��UD��%�pi�`���a03�ٱ�l�_5L�1Go�@s_*��N�G2���y�b]Y�ƈD�~��pѐ<W�֮o�;�t�K��j\ϵ��+/��	� �Blq�{�~�4�UTƆ��V����u��Z;�D�Ư���%����-�[W@�P����"��b� &`�x�p1x��ig�y��n��h�ݱ�(�6��ښ��!Y�\ٱ����|�MN�oSyQ�:�5�
dsv�Ӱ�!�3]��C�H���7�H�C��uX*���)��Z�7Ο]��_\��ʶ�6��w/�W��ѱ����Q��]q�2��>�.��t�w��|	&BAF�J����':*�L��[�(���Ɩ�Vi1@�$у���I����<�r)�d����FܩVtEA����^����Ъ��+@���Ezq8x����;� hPC���ͨ��0`�9MR�WS��+�"�^�T��6�{��1+�#��0f*� S��i����aŋ(�#�UPA���w젡�c6�Uw�l�fvv��5�����*Qw��'2�NV,qG���[ M�B�����|��M!���fz�
�<of��C���]!&����o-�gH��߷�|벳�#j��^j�:�4Vq���?�#{$���u���𑖌���L��@lcIb-� ��r#���!�#�d�i�E��}׶F�s'����⩓}�6tՐ[z��	��$T`h��BѽH����%�,2J��l�z�H#��1R�9t�C�K�M|{w���wBv��ǋE+���"m�]ǩ��/�BMkp��_��mh"D �.?D��@�
��Ed%p1���I��t8J�OkƢJ+LM��V�����@��`xSB] Xc����n�0��!J����TЫk�/�O��v�p�R��i5d1����ƥ��m FV����߲���R�2����L��q�I�v%��t��Z��1# �U}��=����[` �VƧ����|�s��v���$�y�W�'#�L�)-��R�e2'���oO-ᵗL��z�,�8f���Y��X��ytX{�:�2�����\���;��h�t�ƾ��;W�0�o��ZWֵ�.�
`@�ڃ+Eyi��i��T�&bv梦K�}csd�'�FbE�fΞ}oM<K%>�,��+ո{�6eC����a��\��^:zm������et˲��2ö]Fb��#@�%SN���%,_��zu��5�L^�� ���`C���{�.ަ�v�{>��RD�2��n�9jK���va��%I{��n�r������ck�ֻ1K�A3���ځ;���0��L,j���C�:,W:j�}�>גF�+�t�=�d@N�`�`����B�Qk!po-g�,�V�>��6L�
Ԗ.��f��Q��L3Ԛ}��ʶ�>�D�b[̰�,4E�
�mo�NL��/���L)��0��9��d���Z]$���\���IZ�mk
3������(����J�(�S{���}����Q��(B[v�n�؉W�Ј��m�Kr��fؓ7��pq1��	̢
W�r��H8&��'2��%}��������9��� ${�u+� C���O�^'����֛�.�Ǹ�AK�?!ݍRmɄ�Pc��7VYd�����a�̼6����B'M3��z��jW!-�Ҝ��� �A^6��r	�cC1R�9������`�s
^9PV�Xt�=o
�W�_j�~`C T#��F5?���[fz�d��r?H����ˤ�G&$/�N�v�������1qu�edə���T��R�P{ZZ���"��4�a�׆�]��Z[���'�k@�k����$8�rr�p޲�h!�;*�9܂�Ѝ��C��v	w�#)�Mu+1�\9گ�5������5���y�nD�ݽuH�t(�X���d�������t-կ���N��i�2���	U/Ϡ����Э�>�7M��G��-k{����������qZk�O��&�MNkǶ`d�~�]�:ݲ�H;ѩ��)TP�o�+ds���C�sv"���`��&w!+#ԭx'��]*����� ��WgN7�uy�x� �#"\�ǣ$٤��.�T�B1�C�y��!=��a�޶	�d�3UL��\�2$���#����i���ҤL��.�弫�mWY)��������M]w%;�� �	�`�
'/�T�B�[6]/qU ��)�+�/��XVw��s�����qc����|�9x���ƵF�弧�x��椾��7�1{��
0��p�nC҉4ѿ;�2)%�|~��O�؈C�H�`a�R�n8(NI���^H���+>��	���k��zC]��|���z{K੦^�oe�'H1���\��(=BV
<�����(yD��g)my%�gnr!L6�ݽ�r��T�i/k�
T�t&�:Vt��3��R�_שZ�@-��]d�S%��Ջ��_ES������m��c ���p,��c
�3�X�
ʫ����᪀��P���+��ΰ̠��ֲ��ht�.�l��$!oE"�����4������BP����_/(UR�^쇎�c�3Hw�����}|����5��qH�P3��M�Ñ2�����V�X�m<�>��L)���;�C������	��e'�O�\�>Ct�ZP��t]��{��E���W-�8æ�P��ʸ�z�g�H,TH�PQi��E�>1�$�;�|�H�mm���e�@�0(^ռT�g�/��r
|nc%/o��f9�ӳ��?�;�g�KkM3dP��OI$L �hj������>��H��MD� Ά9�p�j�ӗ.��8yF#)`�#_�y��jp%��P�*��-���J3����d�v�ȯ۫��7`�d_��m������1փ��
nSZZH?�~�b�:�k4�>�y`��Ffjc����k�}(��&L��4�]>76�ˤ-L./��"Ӳ�M
.5Δ�≻SI���д�*�O��&��x�UZ�K,����z�\��zIGS�7�y)�+���!G�庯���"�o��#�`��*+&t�:?�e��ڑw�G��h����/P�(���a�Xl�/z�c0�V�����F솣�q�1#7�Y"D�0�>T-3R��'|�\��e�Ż���C��We�b�9k�9��w�Fdao#;U79(\c��>�%e���Mn֘/����ͽ�sCn�w�b��ʪ-��(��A�F���/W��]aX��Y�R2����
���Y���%���q����ȭ<k}����J]%�a�3_"��&!�;�Ŗ��]�A7�묻��<��k��-Ū�0����T��ݖ?�]�b^IL��p�M�_����<;���onpa~�E�ۏ�%�����g�X����>i�B>mf^�I��O�r����R49�U��Y�@Һ+�D���(x�$6�Q�G�􁐾܏GL1��0Qں��.n��wR�G����nw��~����O�S�坏K����}D��[������� ;G���7Ö,�t���=@F�Gt�Z
�<"̓�;�	N�
JTt�1�AV�:J�[]��� ��Fch���]��Hg\DS�|U��}(���?�U��;��t�6\XM��uG!��ZT�όS����E:��)�5W	�������sڗ?ё�ǚՔ�)�,��.[�X��Q�BV��>��ēM�U޻�P O�]��$OR��k�o�\��D�;���9̾a=�|�w�	dp�چ�A.�����@��)��*����U&p'��iE�x٢`r���Z�xD.�z��?$�rh�-�>�be����7$,���'~r�03���Y�G~�4�+	2(*Li�[pl[?������*��
'���Q��|I�:�:�^�8`Ms9�S����Z�$������.�Ej�A��չ�x^oXo���qY��=�^{�����������;��JT:�+iZLN4�Ŵ��(n<����5���6�q'�׃�&�ЫM���T�C$?"�!�+N����q���k=�u�rad�!� 
N>���CDԬ�|%�΅�i/����[��\�1�R�GU��{��u�(�E�5�
�QB����� �|=�m�	��+g�s�e:O'��+M��k�Z���F���Ivd��p���MS��a!�Q��Ȋ~c����Y����U
�~qA�,!��}������L��+����)E�����L�<��4�)��+M'`d(r4P�_L�ҟg`�p���Ëխ�6F|�Xd�2�]��MR���A`d��o�U~�:̉�Y7}t��̃�=�)�.�dn�5 �\I6K\v����!]X�;�9�Mn��mͤ�GHM:P�OE��"Nr`�Ԁ�آ���T��Q�����t7�aJI@>g�͡�0&m���&i�3<��l�u�Bh��+�;5rl�}�]�׷9S!c�
Q�N�Ѧ��q���jp���u֒wml[0�2�HH,�6�,_�����nV�^o���¼N�O��ɍY�4���}v��K��i����9�U؆,��<�:'��aO�l�l��}���xBk�4�� �(�a)�ֱ6e��챊̖�ĵ��6�ڕ�{x+0�M��ʾe5CH1$]lV
�޹"�<H<���?m{H��|�?�/�u@�rx�A����PC|���Z�D��}���O�lm6i�6���b�����7�d����?�Mூ�6M/͊E;��P/@��Q �]�r�-D~��f��gXG�O���j�v�~�/ooJ^:�'�"�'Q����}4��!���s�G�O'R��)f��}��	X��3$�܃WQE��[�������Zs�JZ�Įs�9����Y�9mu�%�OT��z�Z-���-o���atJ�O��p��-*/����;���6Q�h�Bao+o-���4z��g"4\���cm�me�Ns�R�^� Trq��79�y������.>1|?ԲS=BAH��w\Jx%D�;Zi����m։�4C��r5@�<��5�BX(�h����Z��� �n�R��))3������7)BL0�ºˣU�DPՄљj{xgB�R�����'���|{�o�p���X9����Y�%lVn��~�2q��ʣW���V3�h�C�Y�������5P��h���6aȀ:ɀ�1�W�F��u�x���T܁7����^��7uR��]��������)�Z0��C?���B�r,�u_�����x����]��{�2��y���O�.7���E��r?Y	��W����r�0�x�p�p��j�#�a�*���l�ʼʗo�����Mj�"(�{.jE����!�>3M��urX=�zwN:'k�A����kmyA�?�%t�y�qѸ���'�d�d�)V^��nv�6jZ��*q�9E�~;��m��w�'��������Wݑ�:���n�~-P��3�3F��1�1 �&N�D0أ�>^>��;�r)�?8�ĭp��Q��
�۪g�B����>h�8���B��l��9.�?�OĎYn��P�m)��X�L=RB<Km�5�2Y! "�*<�l��pC�Щ6�#R����y��bhq[�Xٝ��� �u��-,�e�+���sb�ƭw�Ve��N��`Wˀ�V�]fL�C��3`KE#6�k��e�T��1�;o*���CC������E��@0xa�K�l��������V6�?-ʃi`�ql����{>t���3ͬ(9�� ]Pj��c{<���k�k�B���OU����� ;���P��_�j�J#����6�m����-�@4Pn��r�Z����+H�?�5����,ߺ��M���k.�X�,�h^���b2�6ʟG�jخ�$2d,J��Ƅ�����
�n�����b�W�.��J�*�ZV�Q���*���(�[d��c���r�qņ�j��A�Fw9L��)'��!�]x�p����XX�(�1)�,ç��tr����7ȷ҇z��NY7�(2i?�f�w���5�I�S�%lɐ���-�<�[`���6HH�tv"���4�|N�~�ر����gW"����� l����"���=�W���H4p���j� ����K^#����o4��,����z�t9�p��t��X��r웙��[XlxVHYEB    6d55    1260TW��[r�ꀐ�q����+�)8��vl���>�a��P;����TpO�rY�&�?�i�L6Pd�+�7ܪܻ��[8�&�6(|~��睖��V��d(̑���HB��~���-��2�֟9�F�=x��,�t�������\���%���z�q,����E��:ѮDX�%���$�T�>��`�2����k"(�i�[�]�vn�[�:H9]�,Lr�޼x�y#O� �OTS{���c`E�	��!�f��A��]��1�� �5�9Y�ஒT���̢�<���=Sa��j�2>ǹ��qB�9~����[fQv�PDJ����O��2���;�Q2�9�6��[��T9|�6F\��_h����	��ح�0l*����1��ї�g�!�O���p���U�FGb��><Ǆ��n 8#)1�!Y~��ةc�:t���p".�_��Y-.�ź_Ɉ��#�{{5UaU'T6@sEMcu2U�PH���E�T�p����+NG�����=��H���a3��QB���#�I��,�ǃ� �]'6��ܡ�.?�0���i���(%Q�.����<X�]��;=���㈨�b3�ca}7{oIQ��<�P��dڠ����ԁY�� E�G����b1�M�Mx�5�|���C�Hc���8U���R��f+l/|U�lAg��A	%'�(hR葮v� ���:ț���*�c�*�`q0�x���afu��Ϣ����l��h�l��B��e�Z��^��AV���l_|�0�NQ��G���Y	��ٻ�#8����3��m헔.Lx��V�lLź��`�؆HJU��X>�oz�,�8Aѵѵ�~�� tx��!�Q�^�֐�z;wG�z�Gz����������Z2�I[}N2�Xܓ��\u��M�����Qi��n�7��t��)V*L�Ŧ����4�̰�� S(�,�Ph0���/h�� ��!0��lֆ0x�>	"�Ȅn�	ѵ��F$�Ol��]���v��c�6���g4�I�NHKo)��w`Y#�>����S!հ�h�/bk8���6�o{0�['��ԭO�{ }�����L�=��,��`��G2_,��c#���z����٪����u$��%*)����� �Cy��c����zO��9xhET�Ĥ�3�|�`�D�\D�wnT��s� ���Q�Յ=�]9'USőZc��"dV>�`y]��ւ6t��*�	4{1���� l�ޜ��N�q6�05U�(-����9\�K�H���T�e�+����JE�O��b��o>��<�-�}T�w���[��s{�� ���R��ԥ��0;��v�s��H�SY:��rg�h�R�G
G�{a�Y��{�^<��w��fP����4+V8�#�P�'1C�S���d룡,��R%x���T*�f*ƹdOd��h�/�b����tN��p-#�1� ��hv�.n�0)�w>@�u3��a̾%�^b�O�H��Q�&�)I{=F���ۜ�T�^���ؿ�d��^e�2ގf#�${��D����n��g��`����������s��6��D��A���	�	BȘ1k���@pᑶ�.��@�<f���q��2������NAu�x_�>���0p����<���>��e�h���]�:n7�<�wvu�%�h�f~�"*AFEB��J����2/4;ns�B_�/���	�O��} �j��\�u��_�&��IU��p�ܧy���:����0�B�[�܌%�=�3k�㇌��r��~���I"�3�H��E�c�Hg�1m��%5\����kZ8�Ʉ�Y�v�Y��ۃ���l:�7��r���a��h�$�`s}�S��)aH�1�Ɵ�o��ܻed ��'3�O޲8I2��� �<k�}�����a���q.F8K->R����1uѕ.í�ԕ�E�~���ms���� cũ�����B���9	�ٮ�c�����z5!�c<����er���t /�l�r1�,}��<@�$!��"G�9��.��F{�zJ,x���c&��A�WlD
KV~Ի�s�a����,6�H��OI��W�����Yߦj�!kP�I��<�<��d3#f��sUw�Qb�~���l� �C
���W�j���͟޼��O�̙��٤�5=R��C?��W�vԧK$�,n�Z�!��)�ϯ�72��V��	���������A*��(	��,c�����$)�y�|5�ېC��\!5��J�E���%��Ӫ��}dmZ�d�?6�AE���9D%^cX�r�s"³��Hr� > �G0�vώw��Mzb2�)Jܗƴr/vC쇊&p!Hjl�Y�2k��p�~�?��F���Y%���Ӗs���^�_�����ms&Up���|e��o=�+��4o�.�UѢF�
L���^�������Y�Y��-r3�Pg[�<G�Frg��x�B����8�>I��ĭX =l�kE�>�	?]��Kgw MZ���=���� q��ⲱ����)��k��d���gO��	;�g����#�5���.����k�mi98�7���l�A�TS�j @]&��G{Hos��G���-����-c��[��vY3�b:�����F#��Aq`/Ÿ3���� �ό���`�k��U-`3rƎU�|d�����tn�L�U���t<JP�Ũ��+���q��ʽ}
bƦ�k�M��ߛ8��:�z5N(�$�{�t��v���X���FQ��=�P@�Nu�"��q��'􊻶R	�{����]�/�/Ҝޢ�`ߜO��qs�!�b���sh��m�u��@;�U~�?���`��]`�e���Ӟs��%��5ůP��k���K��"��)���s��ya�h��~)[z�?��W	W��ϫ{�\۴i\F&��h���pk���0q&]���_$ZN�`IoVI�גRT�qR���Y��BL�9�֧cֽ ����I3�^��'��`�G�n$;�!�S�|5BeBFdE�N���{��.3�#�W�S�a��S}8g�v�'���|a�Q��t�g�!�L��Z_7���[�U��τ%�Xy���W�)��M7�$'�z�τ甕'�]-�y�Z1������)נ�E8~��PM��A���&��{p�C��&�������@wd�j��~R3�@�_���A���q�B�9s+Ifĳ��r̋�)iߐ�4>������p�	g0��Ғ	V'r^l̓ǨD9������˫���h���Rh$��/���������)�S{cD�UCI��P�>s�t���Q��7����p{�4=���ބ�3d,7�힡D���]�����YfB�t�c��ZkOzQ	�ၗ�P~���`��]��5�*�TsB�e�0U�f�MF�:��5q�gT[���H�������|�D�y��V��M�|Jg�0��%�l����h8��6ȕ�e��w����PXݖ͕Q,��W���7�ei=~�����_�LK��u�w�JG�@3�u�~�gˢ̡	/.��-�?�/V�],�� �8C�,l� ���_ΆZ����n(�u��J�P2Zo�x���W��`k�d�թ?Y�X��k��m6�ܞk�8Ae��>��&������b�<2��л��!��S�t�Z�! B}�y��wd��L%�ﱄ3�(���Nv���ﰝ���18+Cl�z��6n��:�m��6�K}r�Ns�^���\���f �|���EFe���a���SpK�sΞ��Y~\h����=��Ag����ӃfG׏�t�=�˜�V�$hG0t_�>�C�~{h�Y�����Z׉H׼6l�d�L��=r�%�|���U�4���+���G­u����ܾ�_ˎ���-�>���,;<�9�:X�[�^E^��QnF�����$�Z�F��2���A��tLL��ȯc!����̖���v�i��Ӹ:@�u�W �l5Li-�|,J7���כ7�f�\Yjf�X�c�B�{q*��,]x��G	CY��v�Vv�Ÿn�����
N3��y+�\ڜ('t�G�|�z� �E�)5Gi�E�֨ʖ�~ %�:�d�ǻߤԎ�^�t2�R�"V	o���S�TQ�M�ǻTeD��Y�`F���؃HT-Wb��'���*�U�q8(�9�	-�e�#��>2!�d�o���*��=2>/j�X�[�3��G����,K���I0�]�>9�[�~�E�e3�0�v�Ȅ�}ix���C�àQ�.��ۭ~�lʒW"�w�W�8j�NT�}���~����O&�{Ǧ����0���JR̚�r���j"�sƖc�E����p�{�
MP��3ՌVLτp`��?�Lk��_cW��~~�( �T�?KKZ�_�F�;�#v)�m�K���r��������k��ьZU��(G^�6U���*��
��_�>�R�L͍C����L��s'M�(^��ˉ�UH���кU;Ч�(����
���B (�m�}OFj焇~JN��Ng,r>�ssT?��
���.M�$��~ñ�+���_5��\�cW��8�����q��M���%�N�̋0��`���6{-��C:�q]�@�H>�Y��