XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v?$�Dp9���p��5��}�����=Sǩ�i��};�hz���X�}˔���ֺٛ��¥v,�����._}�Z�m�H���7Ӫ	/����,M� c�3��t���!`Zyǩ|)�V+���Y�� ��K+�T
����e��f�VK��U�6h�J.�WT�}��ؑ��9_�5s�,+/ڋ�$Oy���i,/�_q��H��q�>�����0����n�~��VH����|��b,J�c�i�8Mx#���%phL-z�N'��+�����T��f�CX��4S���k����PŰB��u=g�����np�`nr���@ݕb林�����ή�tE�ѳ�~]��d ��W`����"�kSބNڎ��검��ŗ�%]��1��jR���L���e;��@(���*M uy���\�xtl�e�j��
K���������g�`D�-����.���j�IĐ-���74&8�'' d����e���qxwj�8��nQ1��~Z�k�T��Gh����{ʮ�y֡��H�=T�Ƃ�ip\wfL�G+-D�Ê{w�7����=x&�"Ob����47�(I���?�^��L�����،�SZ��'����w\��Jvl��A���I�(�%�C:/O��*���@}�bR��d�<uA�^���������y��5O���h}66>$�S����� #������<8;��e�u9?��W��n�v����{S���ϖێΜ�)~�u���ИXlxVHYEB    fa00    2910��)�hr������b��}�[,�N�ø�"�m��þ��J�M�6~��͈�|/W��W�p{�g�V:�у�.L��-��������5H��]�"?e�5쏂�`ֳ�V��nM�%�ӺnCT\�P>+*nN_���!l*��E�bC�{�E�ū+!����c.H�67�͟.�F�e��l��1�k��Ka{ڪ�II�l��^h�
s���k�*�)�nջh6�f���*�bf�hѷ�vM%���O	�nx�����ǌAq|�6�Tj���>�D�َw=��>tK�3��6g���J������py#5����������x8�Z2�q�4Ž��V7�R��[�����z��>G9o:���di\y�4!Z����
B��FI܅q�� t�~	Ϋ��H�<��װ�����@>�k�����ϱkG�Ci�Jߨ���2MnGl��d*[��8]�@HAflB�Y�\���XH��t�Qp8���l3[�}e8��G##.8U��=����_�%��@*e���������`��g�������C3jK��B�ᄑ�=��q��s5�|�P���l�uynw�%��#�Y�8�����kഡ��%P��'̴
��W���{��!`���F�u�~!��ˬIU�ɀl��������G#ʛ���6��N��I�y8�a|)�i�3	�Ș]�0�O�U����|}��V(�C�j��O3�=����mV�	N��I��1(X��w�.i�X|�::�xx��W1
�ѐ��
qeusba|�5���WUq8�V�2Oh���K9C4�g7�8C������B�Gx@��%����*�K']����8Nu�_�k�Qo�V_�1�w�k�i���]���X�d#C�a�ubl�j�rb[�Ju`:S����zǦ��ι�О�.�^N��7��_���k��v�A 2�i&?�%�7����D�Vrb[�]H9$�?�9���Y�.��Uo{���3��￵Ŗ��k6� �^h������Z�BZn���{=���}eC������>(��M��_��ڶDʵ7 @�3X~�甜NK����B����j�FHŋ����(w��A�����EB�6|�8���W ��0>2t���]pϥ0 m����`D
.�G_#>��N��d`ο?���2"��s��L<�>M`��ML��_7k����n�.�������B�C.��� ���o�ȼk��2V.��ߙs�����4� #�I�����$R<©Z�����N4�x(<s7ID�?kā�\�ط5h��ǣ����vS���i�(>�L��b��i�E��r��~���NMO�f��&a�X�I1^����2ȋ1�i�k�uH��"���{~��; &jP��K�xe��\�[����f ��h"-~�iOtIO@�Rwg,�<��/�<�^�����u�:�S��1��K���2�ιA��ǛT���8�Q(g&]�I}e��@^]�y����9�U)���Fɠ!,+�$[Sz��|w��'P�x�l��U���`�f��I�3Y�I��}���N�g���j�$V�Z���ö%�}/q���ZdN�+T�0m#�-���TЅ�j`��2�pѬj��'
�{*�6A�	T#��R0�pҁ���zν[��6�'0�OP_��XZBp���ic�y��� �|�k$�P=d H����#cn1�k9�bM>���8Zo�u�U����u�z�U_#��́(OS�n��߸->3{�b�Gj~�O鹇I�4ֺ|��`\���*�%P�O�q_] Cyc#�jI/ซSՇc:��o��n�����1�X���"-E:���B$G̡y�A$褢?�`�@�0���>�e�����`��[Y%�A�Q�m�5�\���J'�^S��4�	�'x_[!T�:��ᐝ�+L)+]h�r.)GoU�}���"�Ai�=�0p�v<���)��w��m���BQ�A�vk�tǌE��Mk�}�C-�ܑ�s�)&;�Eg��;���������v��_mH��,"�K��N�"c�$�"<�GG��2Z�5���U��8�{	��#S�=S�� e?��z�:�y����E���/�Oؚ�Å��K��V��E�²N(�Li�;&Z��s�L�a�g�by)��V�ǁe��j�<B��5�T�|BTx��?8�}�-��#$t)Ysݙ��N�=ט��41��A�$&*zJ�
�>BhE� �5Ո�Y@�UIpU�p�\�x|D%�u|��4�{T�{���/Ĳ��� ��=��.�2��Q�M�I���c��L��٣B<73� ,z������yg7��_ﴼ0q��''�H��?����@�ݔ3t6cb��V�g$7�b����3 z�T&9�)��4��0:��7QЖ�_�gN�����^Mc�nc�$D��_�5��)H��I�I�����:	� \N� �oo���f�̤ĥ���R��Ӳ�B�CleR��@Q$Y��[k%O��#�P�3��ڰa�ޞT;�[��b��\6��+-YFŚ�TΛ�tFu��u;4��ӿ@�K��D��AkuF��[����9�&K�l�v�;����mKw{.Rt���(����ځB,JԼ�z���0z�	Ւ�5�-Q
9b�57c��ތ9^�(��A��L�ũ���!�c�(�*�9Yk=�GC��8N� �ʹ m6k����)�¬������{C=���4���t��[X�BS
��VB�������?�oz=$u~4Ȝl�#�!�?�]�j	��T��� ��0U+�!����+N��(�.��!>Az6�N�'��3#�Q�R�'C�O���TN/�!�>�{��9 ���4n�l�y��GGEr*=����������.�y��"YfSb��������q ���&���V�!HҖʄ7�Bij�=�k�_�Ğw���@T��-�ge���uw1�z���.��
�����W��4a"���%*��<e<$� r����q���/�*!Ԏ��|��#�73m4Vw?"��!�N�>�d�Y����{�M@I��?��=�R��E�JX�:��R�,����Z�N����\a�Q������u����xA�A?�[�v����z
^�*�j}V�.��]�G�F�çee�i'�f<�1$'qI|)D���I�鷃2���z�	�\h��ɤR8�{��^�_d�ǅ������8�k�7��{�����%8�"�¶��T%��0�ն�W��.2s�Zf�i��7{�*9=����}��L��Y@��CQQhʥ�j�G��l���ʤ��A��1��YM�ʑ�,ʚ\�O.�U
�uW>B ��t�:�yz�r���S�e���]�;��,�}F�Jr��2R^�ϊ���Q/���?�"�C��i�[3i`�����+�Jk���̍�MA���V��o1�D�RGSR#Z��C�H7-�&���5u�t��6x���o�O��O���r���Y�c̹���&��(�����*J���=�.��=1�î�����ޫI��y�O��/|��������N��u�(���Y�q�m,�����GG��3���9�R�J<#�9e�u���޴�Nj�9�ű���C듮 �Li�ՙ���+*�����C�~yVm�"�y�v�T�֔��\���wY������~b%g(K!���.q���4�T�@x�C{M��j3bȷ�ћ����.c��-�#���ÅYf�ܲ�T��\��f΁j@����"��Ĕ��bH�#j�4&����:�ܶl���I�@L��Ĩ(�)�jO�_��^G)h�~&�X'���ᩛjcW��m1�f4}^��v�������y��G�Ɵ�.�y>���@�������U�ϯ[FncPw�P���&֙��E�&]L�;L���r��OS�Y�F�Ѱ���ӑ-&����P��{]d`~��{��!v��qɷK��#�u�F�������V�2�]*u-+��<'P�P�1�i-�����G��}�2���\e�pR7�h�u��u0`��s�;����-	�����:�@5���<� <��4Y�k�r�	(�ܭ��J+���v�i�5��Ѓ￑�!<�	�Ȑ�]"';+	#�I�Q��];��(3�s�ǂxDx���u����!�.W)�*-z�M���_v8]��ʯf~g�>Y��9YX) �6��j��@�	�$x�E�=<����ˍ����A�4�{�j�!�;t�퐗��c�̜p���R�:��o+|��jXz�ݚ�sԒE����/�)�sb�������*h��~�Ue�E�8ēA~�0�[!��(�}�8���mÖ�����%~v�X,.� ��x�f[V��/��H���E�\:��
v�6�b���,�8e��  �!���Y.��.'�1�������aʙ� ?���ΝL
ߴ /�́k;Jk���ѳ���LP�:K������ُ��1<�4��K-���t�YA5�u��8�?���T13e��|5��,�v�>�׌*�����O}q���;�U	�
F�#hƂK�.�=c"B.��Q5&)��}k�܌�Ġ=�?
�e7�"�2��7m��9�X+�z�p���yN�? �;���K��}�������� ���N���X����B���߭��y!\E|�Ƥ�b�(����c}e�(]xI���yL�_�6��Z\q}͝�ϧ]��+���Ւy�8M?�]l��9�ȯ�Z�#��Vi�ٮ��h��a���Ƭ�	uX��������V��Q`�霸��É6B>[2��Rw�֤C�U���F�)K况���hp����Z{�
����1JN�D��LR!�QԜJ��&ԁ��1	�x���5V��i�c�=���s�A Q���7B���b�"?�x��9�}8�c��g�1��"�q	�"K�N�L4��F?��Qќ�����m�amH?O�?s+ĕP�������x��I�A��rSMF��&V	�0��/oZ4^R �?L5O<�Ds���i�(���Y���MӨ��-�����J�1/'� <rM�b)�����`�v:쥆���	j!�%���>ږ�ċ>W�"#�c�'4A6�ԦP���ݲ����\�6�4fR�6��7�|�w�+�=H/�����l�q��j�j5S3dg�E��},�[NU*�뜨G�RPjD�}W�.yK����x#X4��6�4�8P�]�u�� ����E�@��	5<H�ݵ ,Zl��ʤ%Ԟ�h��>���`i�(��9�`���#N/���羾�����p�)m�1��r[�
���.������k����k��b2����jX�v(�/��O�'af9�mm;�:&B��v�MbOg^v\s�<�>,��;�Q��O�K�H� �u�_ǉ�?�!og����.[9T��7�f�I�&����WI����a�g}/ә���]\NA���&�t��G6��="�Κ�9ET������Y_sn-��U����)%݇�:P#����5�z��0�a�?���lV>e>�|�<�%V��q e9�����kKh���4���S8l�����D����{�s}Iv�`���}q&NW�i�wwf��9�VJ�o���ظ�Y5\������)?�J�Q�Ǌ���rb�TW>"w��̂�����<��7Zv�U�QŖ8>�.�K�+^"jOE�I����)����~lq2����%��üZwj@ڗ�F@1� ��2�>�g�T ��3,���ԅ*�C�Ȧ��?qO\�6!�ǆt�|�������X�����-`ӊ~f�Ͱm������)��Ֆ���س��rmB�0t�^��2�dXF`�s�pڎ��'�#[�'��5�$J�mT8�h��ʋؚ��:�Sug.����܋�.����dQ=��cU��;�*�C�Xږ�������E# ���9�z��v�������Ѐr�� ]4��AB�+ ��=�Kr��n.Rf���r4/�������I��4�J���BC��>�wvV"��2��8�-́>�,��߼�z�,ο�0���O�눏�~�"�Nx��G;*˕���-#KeJX؆ݬ~0���~i�o���@W�$8�J�]��"KmZ�q/H{Ub��)��H��N)��f�0����Ժg�Ո���O
u_��j	~���g5=g%1�L�B��d4 ���Ec�2��p��ۀ�dӬQ&�4d=D�7�n C�b��
��KNfV�Dz����g�������g�2'�̸h�i�
�&��ם�j��6�۠�7]�p�Q~�~3��8.��t�k ���Ѽ���\�����s iP�v�a�"a��<j�U~�m�֗��Ue,��F�iNj*�'&|��F��V��瀣�<�@��� -&����9����~i�5���g�F��^�}<�^�<�{v�:��8������ty6�hn�P��B�1�}�������ڠ nAm�F�le�o�k��w��?:��p�y��;+r���:�Fa�B�?���o�w�p_7��M����+�����1~֝�
�HA����}�,`>Ē����#~K:�X��)�z� ��W��\h��EY��A�xY9�K2z�b�$�2wH}�7�����i��#P=��)�ݓ����ɼ����o\��dS#�mu�#�u��Et��'���7
�|��m[�8mOwe��f�$s���T�4oD�~$�05��S�L�fe'�fU��pk�c1���������A�n�
Oopb2	%7�'���<��(��⧳��c�B���J�o����]n)N�ƿ�m�қu[c	����f�[���+$O�/|�� ��� ���q������2�#��ťH�a��	��ws�!�
;J��+s�j���ٍ;����K�}�H�<�+;E�35������`��y�xȁ�@fF�q�$E�z��Dږ1���3�G��h����ψ��[�?��D�{��<�9��aF��<�~���IKڲ�,1�a�ȡ��>�/�*�����n����;.0�1�$ʆ���)@����r��p�NH��F'F̑'�u�������L�f$�Wc��y�t��,����Zۛ�X����Ln�.is3!�YG(��)�-�u)b��WyrY)d
��2l�,�����1�_�B��m�pD��������s�"5���B���B@fݺd<�윧��[�����&�t"UT�М=)��>�R���	�e<6/'��<j�Feq��ьjS���ӳ5�~G�0P�n�����Tڃ`�!�P���ة�B��qQt������W�Q��sL�nT~R)��y�}_"=<e����H�]�',�AL2��yh��`'
"��Yh��tz_��g��K�#\�6���r�V`
���0#F�}+��Ht�Ν+?�n-�L\Za�,O�fI3�P��f�9w<�
�FQ���s��
�!�]g�8�x�R��}����T�1�۔��}�
�;jEd�J{���PҰ�!xQ��&E�Bi�͡h�cZ#>Xf�3*=�?�HS���[�fi����}㒡�VhcʉFs���A�ז�_�TŊ�,v�~��%����>�WT�a��~�)V�|����a\��=�R�=/Y�� Y?:��h�7sF�K��"���к�|�$��wuB�d����/���`�=j�f�U+��;z��é'曝3hlY��|X���;k��_8*�C���;8Վ��~����]BU�ϊ-���B�٘�\<��M��_��&C��{���{gm�ڧ/�\����M��C�g�3�v�F6���#�#��l-��E&:�	J=[�m�\��ʻ���$9��q?X53�#
�-&�ԅ��2]����
���?J����y���+@ѐ�D�9�@�0��:�m����me��.����G�
�`(�l}M~I��"]+���訷vPN�+�����+н�I���V���1���n_��	z)�^��#Z��bj�cX��A�=hB��*[�b���G%|�(���
���<;���x�""����F?��5 �E@�,�pQ��<0���w�a���{��7�� ��BpW����!�Pg����x��~H<{�az��<�	*�S���>`X����5�2%�\�&�\�����6���pfqw݈��y��*Ǟ�Y	q�*f�d$@�Rh��Ed]�������T�;�7t(�����(x5�5A�W��;����腞���F�]\=�w�#�_��P�PgS��a2&��� �����Dn�D�ݍ���X��-��븂�<v�`w<��vPV�·�\�"�ч�Û��g�G~x8���y���E�ǂzZ+Mɩn���������޿���;�p�ʯ�(H�3E�7�M��^���]< d�<����
4���@���W���%I�����³x&��[Ի��)9�It$=�yn� �}�ϒ���ޚ������3?l�����9 $S.��.UവsV[��6s�	c9�-+H���,i�6�Mͣ�S��_d=O]�Jf]l�1�{�<a��FZ~����}�V��>+3��%	����=���~�P ���l�NC��-V'��<(ù�I�.7��jQ\ �4P�����H���(>:>:��M�3�_�"a�r��Sz"���+�e�Ob5֔'u��%��ҕ&�,B:TY3����G��7��#Z��K�
<R��3��E�S�&��x�/r����8m�oؖQz��Jy�o�wY$�j�n{\�%+�n���{���k��5�ǰ<ؖx�`d�+��#�\zM�Il�[8J6�V�=0����O-���������_c�&�}�營+`52FGr&��������2BG�!b݌�:˚�� �����d����i��L#��T����[������,8F�����
հd�2/'����Õ�ڏΫ�D���ۊ�Ew�3{hE
�;�����F;e,�h��]^��r��CC�P��~�_hM���7p�r��~B����b��t�J�x�,�$����1�u~��.����g��q�4Y����G>���bn9�D�#6$�F#^��(���tI|Fklj�G,T=�uײ��M����B�|)���n@݆�ӂZnvA�=�!�����Y���I�!Л�4� �	.cG¡{�f��aS:Z�:�'�*��Ч��cB�b�; ��[-�/:b��D9&t��ˋ���M�X�/��łG�_	��?C��%���dl���J6J}2e��P���ۡ�K}gꉵ�+2���91��{<;����^߼�m'����L�?��GM�%3�_�(����Ιڈ��F9S��a#�Gf����E؍�༶T[�,�r����+h�}��V����}�+�lٮ̔45CG��i`ӓ�3�6�9��;�{�e��v8�c������*��J]������<E_�%�����p��e7���4<�����92
-�.��h
sH��~Wm3���5���Wm(j5_qW@!���`�	�};�v��a�qF��,L.��rxb����tR��-�ѸH�k��E5��P���3���%��y�01Oe�I:s�Th����)[*r�
�U#��w,u]��g ��
*3'��F�� ������m�}�����l��[�B�����5�!� ctT�՘[�g�)���^|�eH��*#�l�b6�'��.��% xDOr�Ep�������l�5�ي?;�{�����3�L�A%�ag�R2(��ޝ,�����
"c��_W���p��e�~�3��
���\�@u!ꬣ>7�67�Di��D�l��P����Պ��b�����A�%��0*��kb���%�z��.���#��,﨨��g��K�&Sd?�j���$�A%h}�@���v!4ă���1<�x+etH�"~PıU�z�܁]�iK����,��o�i����V%%e��NM���PxP�҆(�z�|�D�![G�A.�-Q�h-�zΤy�;H�M��M;�����n��Q�R�w�����i��v@��So�q5:�")w�7����EY�4�����y%Q��|z�%w��P`�U�rsO/8�&n�� cK�?杹^����W��K�0e�[!KS�u&�@�xXe��l^
E�T{�vT��T�	LExs��XX�ϾS�8Wď*yC��q��X��(�4|O~`�����^���0��q�i�G=z~����>�IT�X������������"c����`P����vڵ�5&z�'��H���(y����(j}.�Z�Τ�0&kC�=	OqvA9�<��VUc��jm������#ȼ:=�5vU)�����G<XlxVHYEB    6184     f80%�UEQ)�3�S��IV�Sn4�u��ŰK3C�W�g�jj��-�ƏxY���UD�������3����۲�.fE��:)
�1�
	�pn�nq8��	��#���a{��łv�
-���	?��
9��0\���
Đ��^ ~kZF��"865k�?D)Ox�l�*�a�f�o�Z.�)��yA��	��_Hu�O=��e�"Fz8*> ~�^��D&�J�[%fŹp.w�\�e�]�+��P(�b*c���}@"�=O<'�mD	mƦD�2����'����s��E��'f�&$_��U�s�4V�H�����1K=�& �-��/�az)�!�O>н���6��m/T��k ��檕M7�@�i�g������RW?OM��I�4LA�A��L�)����?���E:�����myxzxz�7h6���d��������ʶ}P�d��k�ӓa0�^W�``'�ϦtU�qT�#�[L��$���e�y߰7[�����ĭ�K(��{#�^F>��<B|��@`�K}��$y�ء�#���)	���q���}ص�C��Hif�+��wMw%�᠖��$WX��D��X�>��6'S�T�Rϊv��ϣ}�,/`��K�F�q�@��]C�����]f�����h2 �Ȟ�8w�L�6�h2�YH����Kު�}�����k��L��;a�6'5{Y3��,a�AŽ~VM�vΚ粍�c��HHqE�!�t��3�p`�>��kַh�:�s�?�E�$6�IGB�^X!�M�p�CP��B�
�$>��E��k N�ڵo��5/�� 5Kd��k���Vv{�Bվ�+'��Ň!�;J��K��cu�/�R)�pS=���џʶ�
�D��h-V"�#�*�~RQ�ܸ��wʜ�7��Ny�VQۛYuY=ؖ\aԈ���|3�E���MR��ŭ�����5�=�%�Tf�N��e��~�O͑��Y�D����v(%H����+t��.�19z��t��9����+�������-U��w�Vi(�$���!It��� @͡�b~�;K��Z����w}�b&��=Sܡ���GW�%Ӽ�R8�a ͪw�/� nm�]%ԭY�{�����b_伇c& _���L/�G�*=C���Y؎9.���/M�	�0"�����X�)yR�6��{�J��@��>'^��ު�	���^�+�W|Y��|�	
ը�r�P�2��QzF��Y{O�#���wj�,*&A��T1�{�}�ι���Ju��Ld�;Z)�R;�e.r�F��W'Ø%��q�»n�����ln �:��==�|�����n��*������+פ��3\�p��)��Ϗb���z������ZPKd�ʹ�����ٹQ(��n�W�~mYQ��<6"?����se�7��Ny~�)x.�g~5�y��
�(��T�]dc���b�м��h�b��e~�?Y�zڨ�^'M�ru8�ɂ�>=x_(u[�푾�)�D&hb,���/?:���?ؘ����6������2 ��#="G J;#�8_������o��8�%[���G7���:�٥�[TU*V�r
̋K�^:������@�{B�o����CL��_D�Q�m,�}��SA1�P�����#Q�Α��ݩ��WA5ò���.��Vrx[���F7�4A�:n��.�D����4��-Н+��_�-	]|�*���B9��-Uw-^����n8���;���ٝgk"�iŲx=z`��oR��}k,V;a����5q ��s��E9^� +�wm���0GO������@�t�79��(����i�:+�Lœ�\E��53V���*G
�n�1�$��b�7Q,�}��R���?-����Zn�#��q8��U�[�KǛ�޷�q���x�;�UB��xb��	�Ċ��ڣ�TI_��z�7���x�Uv��Ū�?�0������g��X����ţ�����ܮ������LIio��ek�	@���6�ɩ�L ���4��	�kl�Bc��Я�5=x�!L,B�'�X�)/2��K�ջ��>$}^�Q�9�j��e9��V#mN悐�Ԗ��6G�Ȣ��[uн�1�nD�,-�	;+ZD���� \������l���j�sf��;x�V�}�K�?5��6TmN곁Y�����G4�/0�W�e����Cv6�+����"������}/�ȡ��Ү@��0㮁Q�;��_TΕy�,�1z���,�?xF�ҕ��i�M��a�	�p��<��mg��_7cq`s�ȟn�m�(㼗�%*�������5���������~9x1����͡]|�EK�@c�C���͗P�*����Y?/N�]�<���5-e�}���q��k���>g�����u��9��z��	�J�����`���n�;g>���%{T}�q�i���H�=TA�)[;W��lOArCDZ�6��!�+���1���S~�Pd�NMKQr 
��H�v�M���k]@��z���\�8Sy�뮻��v�	t5���lծ�g�@Fv�*˿�V����ĪNiC���y���`�Ն!�n��g�P�"�̉i�Y�wk��_t^��݊��D_˒Vl����1��z�t���I��X�〶W{��~a��<A��ߵ>؝��EuI/�'"E�8g�����������'��8����x�E���~; ��OsuV.DC!�M���[����C�|�6j�yW�'��e����Y��\sO�a�W�O�!oA�(l��G��\y��f]=}fGo��L����,�͕FL�BŘ�\��&^��)�p�p�ka�����;+����`�\q��f�>b˟C�`^�����s����
݄�AiH0�(��s��<~�qV���8{U�\�Z��2V�\e�y��`�H=�V�P%��B�rzl��n��X9>���
��f	��K��z��{M���p��c�fb�L1(����yK������9��Y��Z�e�Z*	��'+e�t���:�e���48��(�r9hK��TxG-����֓0���/���+�������A��F�*��Gp(���Po�ƽ��ά�X�	Dt�N�4�껏�i��<��	�FCe�պY����Y��I�9�O���ZK�'JvC�~m]�>�mx=G�"u|����+��YݍQS���2Q;�/��E*+'z��ԨJ�#�v�犐�\aNb!~�N.VedQ"rt��WLk�O��k��12:�i�eJAK����j�Yd+��F��X5��a�nW�%�N_p��F+�T6��SR@�s�ym��'������rb-�"��e�w��l�4�[��D�d����u���xC����<'s3��^%&o{W*�|���$��,Xe�us!���4��L�B5G�^�c>kǳ���*]��c������i��7/2��3�~+r\P
_>o	����I*����� ��,ײ~���?`pg��mb%�Ty���+�vS�`z���Y�Y��v�?!ĩ������X/��,��U��S#C&@P��O,2�{�ע�]�����Ȣ�����I%Q�O��l�4Z����f�|Kj��y�	f�aN%�aa�F	ف_�wyWE̞P��m��Z9 q ��'l[9wР�u�LX܃�x�p٢�𓒜2�Ӕ����X�A-W՗����\�&�����O:T?��,(F,iE�s_^Yڼ�娒ߌ�1�dT����=�W��%�{��.�!���9M�Ƒ��њȞ�Y�|�P:��&�1SL��4��j6����<�չ�1��9�L�F����җgg�~qL�K2K����sE�� �����v�	�Gv
�o8����.��^��iu�I��J!%�9�E�$uq}��2�x���2