XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ƽ��� �:	^x�$n�JU�##ց�MR)o����%��M��ӝ��C��fSc��D�ޥ_oGO�Y+Z���.���614���h44�`����/R.w�;O����jdڍ����NZ��: 9���X=�2/��K���]�Ť;+�mʒ�P����Y�A���"�J��(5 �X���⧻�N��'GZ�n����_�8*@�&+�Ic˘����Ʌ~&��V�L���*B}�@��R�+l�:�.6��j�bM��8\-	
g�b���=b�=��`,�G��r���^.��m��&�aXs9�e�]�,��w�Y�{��2I��ZPޙ:ˁn���e|�Hս�Y�m����7�-�v��; ��홷.��@)�CI%�M�@���B���c.r�R�i������gx�ڍ[؈e������ͺד&5�&�*[wz��0�<�p1l��$��6��Y\�`^�*�en�Ր3k�KM?t�=F��sJST:�$��'j%�6]�3�EK�B%�Í]�U�.Aq�5�2��H�w�K����&G�,M;!�̐�d&�.,7O�
�*�6��n�Գ����*�}�e	�hg�R��yY����Z�+���1�j"�U����U��?A��Z^Z	��[�|���}]�#Q��/Kc�iT�7�ɀY|v,�^�F4�~�C r�q����@n* W�f{�"y+��hpJ'	���_S2�4�`N�n�qD��a����F��D�F�%	�
��p��Al��{Q�:w-rU�XlxVHYEB    5389    11b0���`b:�n-�Sz��W�נ~�'-�2{I���uDd�E�NP[e#���|@Y�O���FH�f����t� ����b�q��~0�c��J=���ݛ�v[�BdТy`z����ɘgƌ��~"�h��W��P� ���褦<B���q��E�߽���d�t�������fۤ�1�m�,���j^�_Fk�-o�e`��Q��n(��w{�S�JG��y����Y�F��jb�x��n�ŬH_DqO5e�_���	��at�&����^��{����^�C2}�őӀ�xb_��iB�s�t�a쩉(Aa����ũ�<**Üx�B'��IyJ�&��.��ڧP��S^^fSLL�\�O�<2�{�S�:�80^Gi��Lpq���Lܮ?�MPYN�܋�Q�����Z�@L��r}�|D������G�M�ʭ��)����̞��F��mpa�T�2�7p��y������+����B:�/Ց��22M}�,���l�-��ݵl>$��h��W7���Aרr݋�#�'.:��-�+�j@Jq�B��M/*R7�P�*_��0c�ʒL�	w�uE|��~ LA:<�<o2�T�{M� C��u�F�����s���Î��6"��Ld���=�s9���{ry�p��R[�
f?�����w�IS0	;T\p��+5|xV�H?�KhdVR�[������@�v�Z�X4M��ڻ��1���ڦ�^W����̳L*rv��3n���@��)�̨�.Z�⺁Pre���Hkݰ��x3qw�S]�{���!���y�-�v� e|�{Q�f�>]t�C���?�jĺ�0?[�r�t�|���B/�H���`T�C>� �f(�9��U�Ōv���#5.��ќ��?	[`q��/�Q��%)�ӟ�^�uIq�t�*\M�Hr"k�h�EY����R�g&�)~w�Ǳ+��21r;S�-�A*	Ύ��.�RC�5��6&�������B�jq���~����0�ө��S�Y�0����,8��9���b\���2��EN�LaH���� e�_毗]��K �Q
U� C	xxM������5�@��I�M����d0�"�"n��.^`b����ݶ@��Eff�B���� ��0
-ȍ.#�Q�l7�|Jq���t-j�Pƪ�ˁo[:���6]4�IX�Gl%� `FL��# 	��IЬV��Z	t� �������p�7��e�Rh�Q��dٻ\*�c,�����V����� ��ˆb���җ�GL+&�3�bJ��:y2342��6��i.~��V����x�{��%��3j�3V�oĒ����~�)�(�]kӀic�ɪD��۽h_��R�2��΢x��7�W����]e�W �9�z���Bw@�d�)�n�	��#d3�y:yd���]�	5��>?1��0D�d�����z�R�ЍX��6�NӪ[�F���J�r���p{�>��6��ͳ[���s��/�*�g�?�p����� ����F�XG�ݓ+\1�>�l�~�sZ�3A����� #��0��E�99M��$�<�o3�Ʊk,>�APr�˗���/#�IM׎]�T�,;T�W��ؒ��/
��ԙ7���g(�1��ǂ`+O�TR�*����N�{��:,Q����m��{t� j���;���L�-@�qv���꘾��1-� �|�2��W�����\��g�^I֒#t��xcG��d[�]�1t��yD'LPE���`�蓪�h���1'(Ϗ��L���*iq�;�.���t�e4-#}맞L�|��ܮ`	I�w��8,i �M�{\�:6�!~�w`�?���?���j� �g���	U�=���εL�?ٌ�/C��U�LT���R�Ǜr�s���%*B��720� 'K��~�\$]?�޽�P�ܢL�ؐ�>W�/fR���sY�Hú���W���0�Bڄ�	�^��Ajs���PÎDaa�7#h�ږ��Wμx��ee��A��v�v�DO�5B�n�C,9���8�q'��vu����у!��F�:?^�-E=86�~#�|��Kz�p����.eGh(���U<�./�fY?���L��`��]q��v�q�z��%{�~8*����ll��DU�>�Vk! |�.�441�܀��i��S�u�}l-%���A®��Bk]�g)���+M";�������պ���E���iLm,���5�W���vm�ks��R���i��jy+�����z�D�#e��{0�$�B��5�Yxq��s��u
-�Asg�L�DN���nk�8.K����2��!���|pa'���@�Y��(��0s�z\��G�P����@�=��W[�3>5f�b;���I�<V�&#�����G��7�Ǟ)f�Qn]���Mf�?�K�ڠ;��sg[�^�v�#��4I�1���u��৻�g�SV�*�t��\��������0��e�V72w�DP�$y�t�q�|��R��Q��ףĕ�S�E���QY�9d������鹚m����������B��x����
��3�Ն�g-��!�8%��_���Xj���7��'3�C�]��uv�@��x��x�YFH�,ZTD>�z�W����$��Z�N��`��Z�A[���4l�X��I<�!JAҍ	]���i�cL�r��q���6'TE�$�'=UM>��ZBv�S?9#��X(�* G�9nLH	��`���6E#E�o�#���J<M��c��OzF��HZ���\�ʐ���2�B"qͤ���tn�'rg��.2��r��bC�U���T�^ו;��� j�#��a.��{.�Ԉ�J3�O���:�G_ޏ�IrX���$<V��M�G�Lus!"u��F�=YP]����ȁm@il�/���%��x�~�?�4{�[�S:{WA�NoK�Wa����vh;nk����k�=����?���e��K]`��B���ҹ�����<v�z�:�}��_�`���6޻�~�>�xq=�h-�@g��kqSw̐ғK�?��5�������)���w40��*X]�-�� 9�L�L�%���uɍ+��}e�c �g��Y�-5�����a��[�Ts�d��� B�d[7ni���_�*��0����w�� ����R�Jj����!R�
a���$҃t����1�C�9�w��W1�q~@`-�^�����	�k�K�����_� 3?&~v�7��4L�Y!'�#��aκ��P�`��{��7���)�lU��wocCL@ݤx��	�gow�V�h?r��:���ȇTEה�F3�)J���#��5�α�C;���ؔ\�K�ý��d0�_G���|���b5�&�R���ez�N�B~�8��3��x������^	6���,�k+�T����"�rs:�}Vҗ����|/�ΐNg|.���^\�OM�*�u!~���fzqMU� ����;��ܰ3勥��59�T�,�Yx�*6����˥�f�&���ſt������۫n���:j}�k��x8�D4Q	iRx�Br�?8���v�^���y)��|�_�e��j2��Kr$w�ZL�J��G{��gx���Q�o�v��"m��%�=�v���2��� �������u��>��n�&c��K�~_@N-�Zf�հQ@���e=�� #���	!9*���r���Jz8����Tl7�q��p��y���/9�u�v^�o>ƅ@jpd3��;2t�X�9�t�ߘ�_��I-9tB2u�=ZJdl?<N���ד��(�أx�SI�3Ve�����T6�\����a z��
Ý1�n�rN��v` ����H�7�g�e<+�^2o��t�ɧ�?8�ԝA,�<��g̒=�D�;=��Ab��ߗNJaMT�������͆��,"�}dN=�``�2n;p�ޮ�E R���4Wb'�by�E��p+�"Ł���7���A~��Ե�!�Pj>	A1�4%k�w-G�2��͕/�ͷ�B��|yJ���n�1%m�����P=�( �6^�d�Q�/��֖t���Vu�f〼�&+{���X��j�^��K8�R�����Yx7}�z}"��=�K*�������5:HMH�H����U�'\50��"r+�&iOG�����{o��-��Ծ`p�C��E(�)fi�t/�BW�ԃk�)�dV��jf{,x�P�L�s��'uP����W�uuR��� �����р���L��itBrO*���'+J�M��5!l�|�;�
�Z�lU�-�c�.�ᱤy(���Cj�x����t����c���8#5�Y'��/'�����z��]L��-�� %�p`J�u���Ԭ�7�6�lȧj��
�sļ�J�����4)$�3��H�ioR�ekt�$C�0L��(�K
�#�ͱ�����fwok��k5���=�9,�rc��:���L��y2��0i	