XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B���\�H�bHx�Y�v��S���#-5b#�b"0�/(􎜓��m�G�`P���#e &��S#/a�{��a<�/W���� �f��xa8��ullr�^a�r1��r��ܜ3��\d/�E~4�un�[�I5d��N�)mpl�hK^^�:z�GM n�[z��ƽ���i'��x�H*�������ԗv� ���7� ��H���Xm�k�.�զ��r)+�ʩ�����z�qQ~hb�ȭ�-�6�I�0������ˢNU"��B�V5���a#�hZ$�&�~�M��vu��X&�\�\[zPn���S����}����\�NQ�!r�o<�ō���A�n~�D�g%W΄��[���J�V�d�Su9E�SC/����?d�zz8���7�t0#|�.�r�l<�Pॱ��*�Ei�䶮���UQm���_�F��@*��v3�xtc����&�=j�W� �W#4�˺�pf��R]����'����`�O�[Ùv?�D�'��Њ�
�?1����jEd���;�I��H�Yt@Q�ku�K�b��m$�օ�4��Ca]���q�* ��M��i0�fF���w.-�M��Gu�IZ]nӟ��o+�?�#\�h�����A�[�� �,V�4d9-�"��;����BT<��	��f�{n*r��� ����D��Ja�^C0�c/E�}��A�����X��'�Bn#�}����<ܓ��M?~ǡ��/80
XlxVHYEB    15bf     890��Z�LC[ȖG�/y�CN0[���\T������zb��<�Ǣ�WW���� Oދ��bt��XiI�춪���a��a���{�X]�+CKŧZ�W��7�gg1�e?	]��9?���$�Z#]��˹׾I�_p���}+�(��
��X��ީ�[����<�Q5=�,�K�=uF�'a�=��//o���~l�d�3��S2*��r�7y��Ӣ��	��������G��Q��z��]&]LX���i���|?�U����$ɷ�*t�e~{1w[�ko�]�nXA_c��u�'o�����k����%���~��3ʧ������;�ߖmG���5ze���y�ɇ�Ir1�e1~�vVg�<g��ĝ0�/��KH�u�� ��h�{�1F.�h�R�v�GXA��qL��\��.��u��_�x�h��xSA�4�G��a�ط�ٞ�e�~������ڬE�V؏�84�����P���-C:��MY��.V֘�WG������94�~�~3܍7Ð|��� �|��� r��r�#o�F8��2۲�).�k�:�|�΍�
,cb�O�<�es<y�gҥI:@du��8���W�� ̪�"�乾j��g1��"Ɗ�e��C��zU���jU]���FDIӮJa5J\�tfc��m�Q �Q�F�rXYjwx}
-A<u��9�}�Ыe(#v�<e%|9�����}��1d�(rIˉU:0y?���[v������WB��QE8�s7�B1I16�9����\�i�
�E�},W����N^��&J]���\�����!Ph�580+�|/��gAw"tu'����D-ͥj��U������/�}3��A޽B��"�űa�9_���XLS[eoI؅���E9�I�=��̕%Rq#e�zx1�,A��
���@z ^���BiH��/z6^�2����à��?�1Gͦч%t�oz����$PC}\������Kt��(�72 ί�@�WSv"�sΦ�c'��\qH@,�]R6��N�T��y�
q��Q�ug��;,���C[%s��zH���ODì;y	
@����@a1Wtm���hbL]$�Q�&ʣa�])����Zt�VU���{9�,�h��j�P����
[d�Ӥ��vǬk2(}� �x�g�叾��u��kрٙh:P��;�=�}��� ��c�P��Z'�rؔc9J��<��%��N����	��u���B}Ѭ��w�0]vH!�����mK��*�߶���y��UY��93��C��I?��9����#AU�v��p�\�;�ō���	�����QA�KШ7��b�;n�{v���HT��x!2�\f_���q�>��ψ��P�E���to���G��۩i�]6{�}p^���mQ�(6^������~�Ł^�󪅖ƣ1�ܑ��_�����a��g�5z��|�eŷ�����62����,.m����݌�P�w�����t^PC�,�\^g�w;k��!�_���N!��4��U�2'E�׉ol�ƪ��KӇ����,h�C/�a�G0)[XӞ���{�3��8�<�Ik�.�.3*)`u��A�Y���a�~ n�R��"�T�d�����i�@���p�{��Jrx`! �QmU�g��?���P��\�d�9�C�a�|ВU(n���ly��?3����zW}��~	H
�x�ތ�~aɬݫ�ۄX�\�fH��m���U�pV�X|J�s�KD��>|���
�I���1�P���W�U���?�,>PMۅ�o�rڷ-��s��x��ӈO�58'�W�RAH�J�l�AV��^C���j@���te���|lE^�x��>�x�#Ox��!�����^'�X!y�밅��T�H�e���ֶgfe�2!X���{�5.����԰���!"ߦ_6A
��4�dY
a=t�����ɑ���V�؂Dy*	�jߠ*?�Ǌ�~���Zڈ�0�ur0��Lt7�c���/ѿ����4�V̜�	�;J�8�Tq����w��By��>�9�P���x��^�����E�uw�?��K0M�"�ꬾ_r4���h}`�`9�u�J�������49-��&zVa	��#������W�/iG���J�����|��#բ8�a�m�