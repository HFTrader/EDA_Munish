XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������3io�Ca�y��C��L�z�WA�o� n�ګ6�2N�Q߅_`��P���%R!��zT~����\���Wl|�.�\�2�,�Q?i���^�*�ϥ���p�|�������D�>2��k����%�t@�LOBm�C�\����5����X'�toz�us�j(�|ǻ���^k}x������z&����ĵJY9j�ha��T-������UT�`���
���9�Ц�P�J��j�P���h��$�O7��Tl��pőV�Ǯ��­�S�1���ށ{�+�� ;C�{����s&���À��u��z����-@�9,�:����� "�GQ�ҌT`�Ζ����
ȥ���k˲�Ԋ�v�(�p��w �U<��Е\�0�*f�E�@W���v/��#�m�E.?'E�iEN:����*����"d>yP��i�I�Wr��%}��&�!��/r���ؒy�k+"QAh�}5�np/����UD�G�&�4��6��C1�S>���g��I��,��l��зw���^T�'sf+!�P�;)o����ca���]2|�<�+��tġf�����P0)�_�zc?�H.��)��d��E�� �4�'��w��j��:&:�Q[�TL���mJ7�2����^M�B�?H��5�E��ܸǚ������� �fVO��Uæ�6w���y�fW)(�k��m��F�!UV���i��#��80ؾ=[���ͤ�sHě�րs@5�XlxVHYEB    33cc     da0��V ��KQ��t�u��N@c4�`��"T�a"��y$��U&7��s��_�xra��"�)�]�vP�=E���Z��*$��(X���8�beeL��o�����q@��Vw܀��4H9���IzP3 �l�Ǔ��9��7��*)�/�����T��+�#���;k���J�?�C<�t�^����t����ɸ�+���D����¨�\��F�$B��ۍʰ����l)&�t�a48��s$' ���ܼ}o��R��m�N�(�O�8��Y:ʆ���I�6IP����>@� l9�i:�@8��F ���!�i-WV��He`,T}�;7�X(�I��8Ŷ�P����=�� �4��}h������9��A��K��Y�H���E��Q{�n�C&��zt�V�/��x*�x�����\���p|�}��{`�s,���S�&w��H�R���։6���	��-u����pі\�Ée�����
����J��$K���!�R����;�R��z�Nv�iid����Ȱ��]! �OD������^��s��[,4�9J�x"o+�ݤy�90�t���l����J�����q�w>���$l�I�֤#p����6��-�
�KUt̉�L,d��=�l��s�'1O��A�F��*�nm*����wh��V�9ڧ��,��%��1;Y�5|h�l���Z�o�be��9�ItdJy�x��1T.���J�}K:��TG������+� o�qԫ�MD5	M6�x��B1:AݚzY��uq�I�v����x+�i��3.~��h��#o���.���ˤבxli�T2&iHyuQGg��	��П�8|K��ނ�w�&��27R�@��h�=�	��tQ$n`�=��߄(mX5�o����ү�1#<cϩ�y֜gd6*����]�����kh�O;8L]]�,^��ʞ��7�����S�����;u�[X���D�tm�N�K����|�zH.\8�ca��Ε=v�#������C_�B�UzH���H�p;�i�X ���=��	2�S�ꇪuzo�/A����~��ݗnZ=�A�����%��-=kb�o�XEs(�W��-�	��&;w.�(�ͬM�Hd�=n�|.O�3��2�N�y��7_N�۟��|��TX�&����Z����������iQ���r�57�8�z �J�^l��]���d�>����X
*1�R�i� ����œ��I�:b9��$<��9me�q[�"\�����,C��E���:=w�\��B�x��)��$4!V��+�N.�������ZurH�!W�qB;���Z�;V?^���V���Y��(���d�l-��DYE|��`K���n����C忿��&s%Q_ ԗ|��]4V��z�ЦV?�J���:�k��E�j?���V�j Z����XJյ��nD�B�<� �yV�q�'��z�!����D(S�ft��T���+��iK�Z�>\hd�j�莘h�M��o��$���{��T#�]��˅�:hH}b2p�ӱ�sq�^ŧ��fR�jʏ�sѴ���5��W��ܽ����sς��}�Oi�Se�x���_�E�4�k�� 1�
E`�P�5 UG]H31W/����'EĴ�!��g���Tl:>��6,���Q��i=x���!��9U�xf����������Kl�6����v�f��Fs���İ4�d���]~<=����J��_��5j+�L>x<��;uн���*Qɵ�U����!������Xv`�u磔�&���SOuw�[� ��+��
�<���N�y U^�p�.pEQ�\��w_�[���a������[��[��'���C!���"���!ka��_Q���9�oPi��L��a�ү٘�>T��
�4咳兑o���z���c6^|�`��E��Z���?в����g����X�o�(�Y)���[&	�j1I��hyqʥZݵ��C�I�g�H��Q��TڮA]�C�P����# ��$q~��.�3M���*N>%[�Mw:|igg�{&g�){�7�L��l���	~(�4C����qZ�9v98沀l7���2��]G�9c�,s�� �xG!��z��,����e�j#h��wGk��7§|����F�'���..d@>rI6F�~�� 6�~Qc>=�jN�{�Fy�$�.}T:�vBL��/+���Z/�L25�4�A�(|6��HY��b6GԚ9���<p)����OYb;�;;�<���2�m}œ�26-�C {R:>��BE��N�E����9xm���^�|�
8�)���:���4��K_�^V� k�Ib�!��CǤE/���P�t�87���:(�������V������҈~X�^̕�̨���dZ]�9$�W��?U0�&���9C����}-�A<��[���D
�n�r�f�H��\�m,t��U�1�_E�UGV�0�>��r���>�xE/?z|g��0Y%:a�t*%���E��B��F#$��Z�3���:����'�(r}>�V	U'-,F��P6��Z����������"V�C9m���{Fg���3�ÅckK�y����44M�����e���B!g�A���B�D4;1�#Ҩ2�;���n�	�F͘J����\m9������
!'�ˇ�Gn�͗�b �URh���&~�@3}�a���zL�'b��K&u�,���C	�6��Ž������X��� FiĄ����v�`�D���ݹ������fh&��Z�Esd�Ed�����R�à���Iz���ZL_�VY*�HY��ಏ��.-�hま7
�`Z�Ј�&֠����Q�0��\n��Z��J2ʉS)�߃�3A��e���<!Cߠ�U8�;i9x0����=���� �-k^|
�����R��	ΨGx~'&#><9vh���@�)M� �d�\u�,�����t���{>��<2L<����π���d^u˱P�$�f�/�	Ӣ5��+}��I�Iܲv��R=�U������i�E-Cs?"�Rl��̣~o��vYw��V��(�A�f8��oD2�Ij^�+f0�ف�kh��rs.>��b Q��M�����^=�����W�E�=մ�#�a��ך����;�n	�1�"�<!��h�k'6�\�G"�:"$[�|�f<��#��$�~�j�������a"��X�	�2��&��1M�ו�u6$�l��:�"��tQ%tBa�֋��������	*=�Y3�
�ǃ�+��b��_�7�Ra"��8>�W^6��s5������	�;U%�Q�`�a6C,��͒H6����դ�S'�\W���$yv�ǉ�D�\���Ɵ	C�BbC��t��b��xRL��
���A>e�y��Q�KU.yG