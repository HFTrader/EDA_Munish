XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��|�[�mm]�O���Ժ��)MJ}�t�#z�W��U+�}�γ���x�=���v��K��n貌eꜧ�㻯`)�2�!8W{ ~e�Q�$��k��X����:�K�� �#���W���Lw���[�MY�� A����I�[�Jq�I�����mi�Q�מ�D(C<dg�ma ��JbW�u=z�3���# ��3��3�y;�di���k�=�l�7��~���J��kW>[��'V�S"�&���ؑ�b���ˑ��
IlpB�? 	כ�v��R�ĺK�	W�ԵU���b^+;�8�C/i�/������{�*lg��(���L�&�8��`�X��{v ���]*qLE�����Î6hQU�<�V���������K`/�N�J��m�d%�n#m��)S�\����c����2��o<�t�5ʵ�ET�FX�JU~�"q��R��d�B7��7=ø�ߧ����#�jGgt�����昗��摷�b�ਃKC�P��%o2o�zpTQdrx�L��{�v�(|���*���q29�@N.�M��lW������Ǜj�R�nZ&�P� �~��Tŉs3ds�m���Ⴃ-{ǖ�4���J��v����"��O�������h��޵� ����{�!���=4�#r�A��țt}������sx�o�١F޷@��KY���%���Ģts�R:E-a<d|�<�F�*�H=�&a)���{��o*����`�ф��4IT?�V~�=��kӼ�	C�=v8XlxVHYEB    15c9     850�����������t�7��Se%�&E�Bfh���C� ��͆�C�w�ߙ��C7+ʔ�F��^Q!#�k{����+�k,�vy^��1l# ���U�p��N VEZeK{�=�>w���0N�W��5�(C��;b���_IOC7�kb�#N�0V<M^�7��"5�cN����A}�l��@�D`Hq��q<���G;R�������:΅`iP�ޖ�l��Ȉ�6�v��������i� 1e;��`ʛw�I�N;c|��BЌ�T�jDqd��7� �M�`��vK�2Ku9�n�C�KcZ r��m�V�uB�]��'��e�V���~��4`����p�[��xOd��t�nD~@���w�~#VW��̇$�Da�~�:�8�\H3���j��}�h<>�I򙔳R*�j����u��(FE��I�~U�r�%��9g@<��%���]P�#Rn�1&A����L*�w%̪B�{Q���=�}b��m����?�����;����Q&�͓���ՠu�x��j���8��d�L���`��Ki��D�&G�q�����sN�{u�rH�jB ��U	�W�E&9�EӤm.Ĩ�]We0�K��ka���4P~,X(>%3� +�[��̈t�E<����7�f����N%Ɨ�ֶ�
�m:����7�����a�
��S%����{��F��/�����z��yCyҘ�(m/�i�j�re�����DME�6S]�"�C�V�Ks[v����z��|ZF�9����#�_�Vb#I �pE�5f��L�A���}mJX}��W>4�<Ь"�T�E�q��4^/!xGA6:��I�<H��ѥ$��,bP�A~��]�y9����+��䝹5Y��a4�oQn���I�x%]S���1�x����ٰ��>H�z�ʚ�7���	��*qy�d�w���u���6�vȑs���m �$�f{h�1�ƍ��֛X��(��߃�r�i�
3D�p�
�)���_���0a)�9�V�>,p�t��~�G�����4w�r3+��I�؁S&n�ƆK[#��E��ʍ�+�wǆ�3Lֺ���? }#�ˀ�- ׁ)�q�HX�?�z�q/[[�^�?G�#uy���]ۛBv�ހ����4�k��V.24z?���6������RIu�gO�Z8�bS��g�19(Hs�D��ŤB	u8@L�i�>&�(�N������Н���ld?��7��F����e��:vA5q�/�[��&v��.��	�S��i��@���_3(F��׾}}�� �3�.^Yo� �1����Χ���g�Fcy���y�*`/�#����ڼ�Iۮ�ٔ���ԅ4�9~�=g�T����-l�߸��fjE�ZH���e��{�:���9@0s,�sAn/����yj&��T<]���.c�'����웴��9������=!��<b=�%m�:�`���}���p�(��ʔ��"=�"���XV�J`0-p�2�� 0��~���V�M�R�H =p�@���J��q�B��=�4��h�k�Z"e��ܴAu��H�r@!L༘��+�ĕH&+����ȱ�vp�|tѢ uF����*?1f'p[��;���^�SK��	��)���
-������3���U�wQ�s:���͌)��^�*�f̆�'R�p�I��-<Mfo���Y�'�vy��oV��v"��=��߽hD��*l��d������OEH�n���Wmf(h�]��������b��U�ـn�~�mf�����Y#�u+�=������A���%�O�o�KEF�f2��y#�Q�h���iJvB�8Jx>ը���
�:�����ʲw����ҕ�K����ڃ8;���1��?�׬}��&�l���l1j��kKt�>��t�,~j j,��n(7��I�����WbH_fC�;t,{c�Z�L������cN�(ݯh��<��
�����EG3n&�3�-��O��o��N�׎$c_�X�eCؑ��1�5>�5��:���]�=ed�/C�;a��t�+��!Eo��%��*�OT6+����Z���N�tG'9|����~G�Ւ����