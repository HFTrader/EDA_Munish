XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�`ˠ�Q���9�����:�m�Y������ R��mz�wai�(��bA�>z�|�s��_�:�ˬ�-@/Uݔ{a��GwN�8@*�-8: h��,��~j�t;��1-�����f�U48��,�&g�?ZB�P�4�h��|}:`+�[Tغb��Yn���M�8x0ת��F�����|{����SO�u@r����J4X$���r���o=��I����{$*�6�qP,&S3ug�m*�?h7?;�4j>������_[d~���0#kh�\i����)_�y�Ж"_�Fx�0�NP[O�����?�;�E�.]��2.vg, ��A�?��	Rp
n��ųX�k�Z�+�PU"���l6D8�zZ�Ϝ�Un�2�!08W ��&$E�9�����@�28��I��s1�Ɲn��T�?"-�x�z�B�ϯw�(O}�뎅�$��Zw��I�h�E�tKBm#oq}��/&�WEi��&�������-i6
`zlH�Dn�*a,z��r����S��d�~�$n�^��y��i���C��Yn>xDq��"�$#��n����z�\� �nT� -t��N�Z���/Y<��Q���*=c�>C|Ϫɗ�	j�G��t��1�"�$��8P�n��ǛҤ֕M���ܮ|צgIxq�;ǳ�A����uRF^'3�g�]�?#����w�s׳*������[3b����&`��g 1�[���z��S������v������)+�ֹT�|XkXlxVHYEB    63ec    17e0��hDY�	q*.�!𯮎s��P_C1�3��ݚ�|=���\��$�^E�@��F����H�;O�xe6�~��,Yr!6�`(9L�a��n<�^;-�����
��M�����lQ����u)��>{K�W�R��S�Kᦄ"gh�
�����Z�i�VodB��O��D�\|��)���⨉�ޤ[�W��RVm�M@���.ep�n���=�,��5.65�/�yFC3C��VL.��k�-��2�5)�5����hh����;��A`'󒄘�e&F>&9�57Tpޭ}�������ӳ��^��@����m�7��7�4brN�!��gO�'[K����BBo�Z����S��K�*�0Pr�1�QD���m"��BK1�2��?��*���ap+A��lF��e"�=�<@�S ��'w��+1�T��
ޜ|V,}�v�&)��%�c&�H�ߚ6_�{Ǿ@j2u����<i[1�sv-��i�`�^ϯ+`�Կ�z�����)�/�|U��}J�"�?*k��3�w�Vբ��eԷ_�2�>φ�3��sw�s�N�p6�o��&�`�J��[4:�Rd�y�O$�2	hON
�U{0��%������1����j���%tp��	�-����8����#���^��;5��]F�C���3`���PK�����8�9ЬI��]��EC#9ֱ-�^bK��N�?ӝ���8+�۩_5����0 b�v6��z�d$n�ۋ�m���
};�Q���9I@{A�FZ �d�SL�����y-wT�IAV�d��v+^��1�V��i�4De6w�t	D�D��E��h�s��P'�!ѫQ6�)��=܅>Be��S��v{E4IU�$|�4\�:��	'>]`���[��a�RM������L�X��`dTE!��p9)����*^�������ZZ
�w�Z��Dj:��K�����	��.={��rm�3F�ɘ̤���0�*I�BRϛ��d1'�0ۄ�8qk}����OJ��w~R����C$@��Zu�2�7*�A2��"��	��QX|�j��~�AB��|To��p�t��7�)(���|A�ν�3���]?�6��@A��P��!H#G' ���v�ܴɇ!���!m�F�g���b��L%`1�h�$�#U��&�'o�o��ЦfƧ.����U��o�x�n���b�MI���
�3���~���$��l:�j������:��%�\�Ce:���`�mº{fA3G�;Ԉ������k<a��.D��#��w�%W��J�d�'+��r�~F��tjy�=��8	JNlX���l�	���{߲���$mn)kDD(�EZ��I �"�>�'4}ϋ�p�ǿ�%�WRA�&�j:���V��5w��|Y0��X��K�i�>s3rږh��辨AA+���i{�<�������O�/l�(YV�B��XB�a���|�uD�<q��h4/[,�\�n�^PC�B���B�㦊��_�h%��F�F��*���γ�rrBl%�sS�0;����E�5~|�Um~4�!�ڽů�G�<���#U�[���<)�0��+����=�`D**|�j���!_A�Ɉ�s��|��Pi�s&�����+u�4�\�-�3d=�=���3���fZְ+���a�~<��r;~��k�� -��Ν�D�jha�����1dH���"�����b��CP�Lz_�=�og�M��VՉ�j���~�w�LA7����Z77��\޵[���d��;�C����8~8��:R�&�U2!"�s*|�Mc0㋬O}��[io�_
���"�̉�}hG�Q�����v[�J�%�$v ����'W?{�>ʸ���jF�������.p?�%��\hq�\|ʔ���kB�=}	J�!���=���f�z�O��v�*è!0F��,�M���L�m���PA�X���1��1 ��N�ń�����^ ��:�BP�r�0�膖�,������Mӱ������ё���^�8��J�`Z�U��8�!|�f#vy�>k�-jB1�fj�0�+���W�Cb��ؼ�����Mw�vA��	��-N���? �ĩ��E�x�����׹*	kwБ�����'����������ٛ�7��*��|@���bN�H����C'z���ɡ�Ն��,�P���S��K�W`�$�s������80�j�b�5��Y��_	�/�ļ�����c��_���Y��#�Dy��|���r��ߚ�b;M����[*�]�Jr���4x�5�~:%3��*����S_M�.��D=��$���5Z6�iA����ic�im6pW� ]��/(�M�WS ��jв�2���(P�XMw삝	�q]�p&;�����ӽ6?�Xcn�v�7�\!E�I�(��ͺ"��
�]R i�#�Z�9�k��#\	|�u"��H��H+5�|�F�����bJ��D������p��JGd�Q�A��]GO�����l�zf��:C<f5��TÎ���ே������r���h�0j��A3�����ET�@�`A$�] ����s�3F*�=��ۨ1~y�6�'�.�i&릇���^H{~I⽡��<$E� �}5휪\�z��!-��}�����X����A;�R�P>F�+��W�e����_�7q�L�;��l_�K�3	��)��ʚ�ԈN:1��@C2|���AT�P�/��~Jr7�4ks� �2b��,!H�Sv(s)���1?��>-�ާ:t;��t:��s~~���w��{P��fi��Y:O��Z�-���Ϫ��jL�2u�%�q�����3���P#�(Oȝ�by�*L�a�VI�n��+�1	C��K�=N�����D���3�_>Jd���]%/��PI�%�K���[�zu\4���AWA�Gj�G9/A�c�gGd��2�O:�|��č��M������0���5Z�~������a�n��L����`��H��p����2��g���?�[1�e�1�O ��%$���e>�O���ے�=���T��؅�p|n����!\< vZw�Wc-ϐX�l�����?�g'�k����Ut�n�Y~���XO������ ڳ�箝$��v�>��� b�p�/"P�B� �S/B)�Z�N����{������~WSI�8x�N9��͡2n�����c���,Ȕm���d>w�˄h��SZ�����֐�c��c��x� ���8Y �n��
|$�XٕY8r]��e�<�n$L���_�c��+�X��'��i�������e��Q"�:�C[�V5u�1��>�4��}.(�-���>�.��-M� 9�3��\��v�"�N�G��dE���r���	=c����;�$�m-i}v��Tؽ���嚱��A5�Pi=HL��5�'(��E��1�l�o��e�1[bUu���>���1`������l_:)@�n�o�������a$��Yj89.�R2(�vf��)��L�3�M�&��G� �WB2s^OҖh��N������ zч�mX���g�\��3��\}�}��K��4*l<�m+|,I�s�)���'�b �^"�B#����R--zJ7:�S�4����]	3k��N��;kt�E!D0-Q6S

�]�h\�a�'�E钧3��7`�۴M��:���:{]F�@���F�E��eĦ��\D�Xe�hd��*�s��"Ԥ
eyh��|V��O�}�ʀS^�]�gF@d��L@X�ju���O��,��<j�i���1��J�=^��畐A9��~
V�����>C���>0�A��������X}��ʩ�D�����J��lb�����fc�6�������E�7q=��F(&�a4��{�0�`ÌV��v�)�{Txk���%�9I��i��{��	���L�5�@��ʕ h���`�4�Є�+���&�V|ߥ�R�_0�Wme҉�(��,�[�:��9�7���2��	S	�Ai�|�~�����
�����wx�2���e�림NV�c�7��n �ťY�:��vIV���C�"V�-|Ԃ�pr�&���/4
���y�Eh0L⃩/��
��I��15��Jw��cq����?��M���W&��H��^�M _Xr�cA�>x��R�;��0L�)ֺ��7͑�
���1�
͎=�{ٶ��`�gcW� )�ރ�Wqڜ3u��"2�/���ë�����y#�w/�vi���h?�,�̬0���-�~���"E�HB�4v�XE�~8�O��h�2����]����3��'`�h�Z���3�|���&��J��b�*,{��&A���V6��!�-`x�Q�Չ������K��=kf��N�n+��Qa�����P�&Ň$��y�i�_ʴ�S��{�[ c#�oK�z>x�/D�A�ᛗ
���}n�S
����w�����+f���,D�W���c%�?��֔b�8G��{2���^�A��aMJ(�xg���e���U�듚:����rpK҉� �vq��>6��o�pg@8t�|�vp�z��s<�Y��Y��-��^�k��.�ωa%�쇦7m-�zm��P[��n`�54��R0�h�0M��f�6N�C&v\i�	s���GGM89说�ͫ�Ԓ��,.��T�eG�F�c���?���*�����_���t�Ww�(��7D�-���"ZN�{{d��ӕP*FKL���S�j��_��ݔ�ڔ:R|ya���Iǀz���f�[mB�a������ζ����yl,wؘ��ܑ �e/��x�W]y86N|�O˅�	�0�|`���9�R6��=���W1""k�zx��_�Q�C���2�1gn)�h���9B���q�w���v�T\q+�mZȳ!0%��Bf,��=���Z�}��:��Ԙ����P5���V,Х�H�Vjt������*Au�쾄�#��L`����,֞U*�:Ψ��Q��x�D]��H�߳�z����*3 e1�񁻐h�`D� /��H�g�p�a?����۱���B���*��LZ3q��i�%R�c�T���"X$��m��՜��������bY�@�|�F�����y�8d�_���F!`�Z�E�[���0��B:��$����v�T�h"����h2�7{� �ٙO����iq��t���I��;���? =�u�~���Oh	��h���D��AFRh=�#{p,A�j��;	>��4d�_)��7���IE��x��,�����
<�)�˓b��2�pi�����1��O�	���Uj=�֞Q�#@�$f?��;���)����t�^n�w��]Z�����?lhDab=4�!V�̋�I��h�b���3�H�����Q��ó�;ǵ�a�,C��B��{�HҎ��ob6�S�0�YＺǼ�C۲y���i2�C�J��=��I�����v�:�c}'mÊ���?��d7 �F�԰'#��ޕ��H}�,��:�q�x̹�����{ܓ��FsZ��Бk��+��R���􅄯rI~� ����I|�n���K�uPZ�_l!���)|S��"�z��M�3Kc"\3�6=���n�؇���2���+�h�]�海�l�
�����bĿ����k�}
D�X&{�?3�N��W�7�E^�[�\�I�G7��l�] �_�R����8�ڱ�o�)��Uz9�0���J�HK�;�]f�R�1�I��hw�N�Y�{sx
�S#������@t�S"��.]������q��|����g��<�5�lc���#����mp��Q�eMi��[g��o����c�W���l�2�@���B��|��%Y�TT~��V�^(� ��@�;��p�oB�d<���u�6�1J?��4B���-j׼���V�AkM�To��2�f���̗\�JJ����g0@_�;�Q������������#�D���?X�Ц�f2���_�������qD3���?�'軩�1�큫�O�2ȇ,HM���8��tқ�