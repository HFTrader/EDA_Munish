XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��GO<��Т�E� ��ؤ���	L��׶���"A���[l�)��!���.ԯ���P�9�Q�v�����v���!JhƘ�g���a��m���pOgK���E��a��Q�Q�&��#W��x��׎�Z���W�z�;5�xAw�}�n��;}L`
d��d>���(�Ɲ �m�Ž�d�0Ի�!�d�^̕���+1-	������s�!�gE�Q����Q{Ƽ|%f��/��u�3X^r�Ǳ�zx�o��u٥��F�3m/iJ5䢒��q_����K�`�pe{qK֪��)�baT0�/�?\��Hh�,���oFLC~ۘ�d�e��pF'��v����S�be�w�%�;XU�_𥙻8���+�TU��9܀(�g����r�Ud�����@X���hV�z�L�e�����h;Ԝ�#5�~W����ݎ��T���D�������V�8u:�
u��j�ʭԔV�(��FG7���.I��[qn�mC�$_Ǣ�ӄp+�~���٬���x��������#��V�|�-n�=-(֧��$��^&&�;z"<?�ˌN�,T+��k������j$�Q.�1
�y�n��cH�ɠ|���$Z���u5y�5փ�*C��K,�;�-��<�������������pke$*^����OČ |�)tsj���Z�h]��O��_YW�@(��;�������!����Hqp�ŏ��c����S�~���p������6GXlxVHYEB    507a     f30���
�I�����G��i�%��`S��2_�`&��c?yz�Aw��=�*F�'�!�˻��G~�d_������;�i D��aI�<�#��~��,EK����;��������o.(y@\�������Z �'7�ٱg	<a�r\ɜBl6�3}s ��E���[l��L�3�=�&��v��X�{�%w��?-�3B��2��qA��O��v��u[�E�4N�UQ_z��j݈`��ap�˝I���A?��/_`fw�e�%F��m�� ����9%5=���!�f��/�8�s)\ÎJq�4[�'O5�ԁ�(�%��k�2�qp�}8��u ec�CmW�	����T�p���CF)��j�x�I�f+%,( (��^S?��x/����9�rՙ��ĩ4N��1�E�U�L��hO\NU���[	��;�$�F�W��=VB6�����2H�_�l�G9�L긽v�nm=���,"��mO��&+��b"y��lr�H�n�O�}'�>[p+�m�\���q���fi��г���Y��)|,����+������Ԧv}W��S*�&�+K��kzf���9�Ʀ���X�}�P��A$_��I� �KH������2���ԧ�"^�I/�=�m.�ۍ	aOΗ�}.f����$�"�#˔��U�q}f�/���C�9`˄�R�^	�^��EȆL���8��}H�@�2��U;�ɴ��؟?}�j�i��j�.g�`��}�T{�E��i)\=mwI�D^��c��@&� h�X��C�*�u�*!���i8[N�i�P�C��I!rO#�N�^�Q�4V��Y4G���e}�)5<�'9� ��^nB�H/a��u�x��q~��>�w\3w���KU����cC*n�27�����t��I����FF��%��Q��y�
0����9��f�8Z1Xr$��3�΍��:����%[A9>�m�us�N'����~����_�:��ĥa���e�Ɍ�%�Q?��K��e�6��41��po�0�`��콻���0q��^�id�;u��8�,��VG��ϭ/Y�ӋP9vػ�ռi��ziu������X�϶�9��hF�\`r���W��`WՉ�ys����Ն@����a��<���Δ0C��j.xN�C�����X>�ݥ+5��������1eI]ރ�}F�����O����x;�i��s�l+�Q�S1�yO�@g��k��d��������)�m�,�#E[i��~Pg�a��k�o�9`�����Gf����O�(B�st���$���;��8��^mq�!� W2��h_��+�Y��
߲�cg�l,)��zc�g	�����}���~}���.]]tYd�<��{�H���Ԕ�S�I��n��!�'�IF�`7�jY��(��Yс���C�g,�U7ի�i�>x"t��f����wKʩ	2��n]��T!RWi="f����?��mC�.Ң*G;g����x`�)�Km��i�ǁxK�o��e��Io�/PK���x��� r]I�`5
�ۥr+x&�wHl��ߕ�U��,^'v4a�w���9PQ�oݯ��Ҵ`���s)3���I%x"�{��+򵂊q�O��'��UUv��Y8��y��/��RdI��A&n�h��n�w���u�q0T��|}� '���U�يN	��Z����r�k
���(qס30��GS�e��0K|6�s��R��P?��Y9mbwj!�-;�y�#a;�Q�D�����ߵ`R}>�h� g��VΙ�X�$���ؕ*��^15��/f{s�̋�vg�:�e��`�Gw��>�Y������%�M��F��"Ƿ�{n�7�v��\��s��(A�eXRMm<����睼��:+������ۋT�K��C������f�e�;�,�r����2����,H�:1gS�Irme�UT�/.u�h,z��r�DG��b#kTs�&}��ss���Qt8J��]�ԟ������f'�|6�m��p�� $�r�E���$]+�r�~-�vS�p�e5֛ahXU���χ�1(�â+4dKd����O�����r~�EB�<U�w��.&"f���Ft��F�W9��c��T�{6�� 7L����W�!]�<�؊�k`j�a���nfB���6*U��F4J�|�㰌��1,YN��ߡSK 0{��!��4t�$��X^�z�;�d�|��X�����j�{wr�L����U���O�'�y���/��Y���r#jG)��A��=>J��|���
	O/��bw4N�ӡ�^���Õ�SymX���O_d���rB����7�y�o�}c�z���=�^_�I��g�-���ם�?
�0D�}2��2��Y��h����c*Wso6�r~�`�1r(�%�I�XtxG����ᓑ��f� ���C���B��Y�D6!�&��I�w����dTf��2Dh��D��L�����0��!W(4��;,�^��{��4���m}p�7�9�701$8��=��$���z����O®��� ��|���Oy��׶uD���we�����l2ZNt^k1ZԱG��9��]z�oJ'��&(�u]���[����-�ԣ����V�gl�^�n&*!(h����e8�
�K��(��&|���=�W�^�]�ٸ>^X�B������W.��ٙ�0�|��p��/`m���6�[�'9}���`�/������������6�6�4�z]�@ֿG0�MXDa�zr]=�ДtC�2��6�A�;�Į+��m)<{>!|>J�\Y��1��yx�O\����f�1�C2��ɩ���*>v�I1����0k�1cCCj�TH�M5(�w�#@1�?;�w��5�l,��
��V���}�R��~9�|��\�����2�����������Ũo�a�51�'#G)��}��i6��\�����aYx����p�'n>4�<$%7_k2���nFz��O��Wț����f�I�[x�m�t�;kV.Ǵbm��v2�<� 6�� ��3A��u��z�&���ߦEZO��B5$�ǔv��i�V9Md,qd;�w=���s�	ŶtF"�·������`��	�ޫ�R�uu�Z
��2髯[(����׀�f�2�w��=�x�}(�����q��R�����_��7`ls���.GǔM�U�\}(�.�E�kZ3*�jԠ��6�M��#_�`��ilW���u��hi�Ä	�Ir>���'�5��.�J�b]�q"L<���w��_���`B5sn��r���<�39��g��o|�ޥk�x���"ճ���H1���IӞ���G&��g��Iˏ���F#����ɒ���" H�����]���;�
/�:�P�#4�p4�&��)��b��ݶC���u ;��b.�Q>��L�fr���N]y��[���*s!��z&)�q@ϣy����m��ҳ]�+Q�������YP�x�����p�K7�~<XL��V��Ǐ���	��k,�̛�����6U�y:+^��\9䈡�[�M![tu6�f�$�	�k�tMG���4���V�U�f݃��7�_��d��.r�Q(�ZKOKs�}v�),cy��`go��6��E��`�����f��*�\�[��P�ak���Su�J�
�Fu���ă
:�;s�_(Q���X^
�K�op}:咔���e� �&!�����|6k�-��>����Yp��A�i��>�|����'��JW��[��E�q��yQ-FRAS��R#&�:��AaK��C�`�;�B�w�p|i��o5ymvc4Ȃ�\ֈ0^