XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5C�<F�XrU���9���t��Ԋx���ڝ;��V�L���*�L?k�)4Z4��,������H,�owT�|I�Z�d+��y��j��d5R�+���k :������V����"\��B=p6x-A�8����f��k+� �Ե�ԝ��h��_h|AՏxE.�B8o�	��~�p�~RNWǆ�=�E�v��$��W������ԛc*�$Hl�`[�a�rR��cs�F�_s�S._c;�]���yP�����#0K� �1v�z��ϋn���b>�)3-X������J;f"?�+�΃pA����aRCV��4�߱"�.Py���r�D�Q�eP������X�E�0�����Im�?|��>-o�61#�ob�A�{�g�M���&�ˮ��L�L)6�y�&�o� �Q���#X�'*�;ۻbd,av�OA�0�s!`ߧЃ�%�\OInu_y�iO'a�I�6{+�oͰ�λ�贋�O{�GEQM-�c;��`a����x{4(�чXav�,/�S���LR�J�.��}�._��A%G� ���B�b&�����rGh��y��O����@kD[��v5(�9蚵��OD��ݬ/�؃F��2p�����v�>��=��Y<�o-���#�)�����_�K�KX[Y���P3��9�HbY�e���p/}��f�C��o�}�����v�����سs��Z4d�)�Q߁r p�$��?�6���\�0�{���#�~������|-̏�Sb*>XlxVHYEB    893b    1e30�^&�K��;�	<L���s��li�K���.�5�g5���l�D��L���S%�?:A�Y�����I������p����RIa����嶚�:��8���������d5�<��Y��Ͽx��p�|�%���yA+#�%D��c�Ms��R�HsT=��O[��ľk���/n~�d�X�Qr���a�.��٢�l���1(30_���6���D�����h�{uz���'���O+�*km�)���"^�C�\pIt����m#�.�E���T���}G*�bb�/t l�/&��9P��J�Ľ�یb���%����DRiݨ����-~�袠��^���S0j阨
���%��͎�a^z&���墎�%���1,�0K"XM-}�`A��:���;��u]�i�;�'�T��� �r`�ےiW��r>���� �~��xl�`�|�5\n��;��;�cG/�ehJy��8"p�J�Ӣ+�D�0�Ȑ�D��]NT�/Hj�ɑ�����yh��Y�-r�G0){����D�UDݾ�m�l�,t����pH�<�;��K�6#�Q�ڙ�k�܉?�|��7�7�0�q}����Dp��O��3K�[A8aIC����p~I'!w��6 �%��+`�i��,7'���N��med��-h��r��ʅ�׮��h�\���,�Hʄ���Ϲ���:aGs�bI�=S:��;x��&E��3�`~ȩ���.X��U<#8B�ٟXt9/wʪ��7Z�+�����x֩n㣔�߼��c��SZ;��f�c�y���� ����r�O�!��e����h.�4E ��&�R�����uNd��+�t
����0錾�U��b�[��g�J.D�e̯�(H����m�QP�v_54��}HA,�� rk�&�x[�)�~�y���!��40]��6[#V-�C#Mt�u��Rj�F��7V�ǖ�4�H� ��j�^��k�ۂˬ�x-<)�^ĳo�ecFW���12b^�3�9�2A5��
�sd}����"Ӻ�S�=�@uy�6��r&P��t�k�e�j���p��Q�S)����1�/���b�gЫ'���R�C?��G�x�������.\��?�d���#���U����?�4�.]�G��7���H�_��N���,n�|�����ŉ��%�3 ���c�ވ}jx�Sa�$I��B���3��\�q#Ï���T��g�1!M8p�a��,�TM���Հ)D��t��S܂:�`u�,�^���'����bգ�|]]�78ݎ���ӿ-���bM�S�d��/@��kܟ�N\W=��p:H�73�q�w����*@���ť|��raJ4?O�2��9T���y�w�
i^)��w�eV��8-'+H�J��$���r�c'0�@ǈ����cv%�.o�L�!?p\�K5a)�H"��lb�۠/m^f��0����]V�S�T�s��i�*��N��X4$c,y���Fr��#���k
�[�#�z;yy���J5c/��M����}S�T�V�u�}�z*ss:ݸ�!;�( �G�T��.;�p_}Q��������Hp}<�O�=���I�9�1c4��;�� �tV(� E�_�q`�W��V��c�Q�"?�I*�<w�W��% �#��S ҋ�B��R�є|�N'�"g�����K�;Us�kȁ�tg�R�N�I�w�
�<-y_m�Gw\n��_���u��XC�|r��N6�~P�}%Q�Π��'+�����l�m��	M����BZ~L\��H��l�H#j�k�E��/��}B��(%~��w=�M_�(�.vVY��;+�+إP[IV�|'�<�*���X|'�p��I����(蒇��=w�j�q=����v'��3�S�>��Q�� TNV��;�����&L���������z�<U��挘$(��9�e���oLb5]���B]�!\�Ys(�ȿ��)8�	Qmo;{����|?�SV�����M�+?������D)Kֵ�j�ڻŇ����ѫ�oW�ӈ�N�<>���;�b�ڼ������D�ݶ�9��}z6��{��� hR,E��h�����]:l���
�[O�y����U!�T�1�Ňn_��۔�#Jڽ�NZF߱	?�X�Ӆ�b�խap�s�8�F�TB�5�é��{�_Z;t���dpR�������S{b�9beUm�Ȓ?xā��b�<W2��#:����T2�z��:ߏU&'bFT�mԌ����.l���/��TqcMOoy�[�W��iqߩ�܆i%�"���5��E5�T�P?�c��
��cc8�H���[�!�xVt�12��\���(�32[���q��jd=���}e���d@�8:l�"A���N����HG׉��7�q�zj�:�ܲJxs	'З�&[3����|�N�K�֥%�ޞ��f��Ý�[�_h^V8��EC�����5 �"���
�a�����`[��ikz�59��^�f}/_�A�t�k����q�m��������v���V/FK<&��?=k�j+7У#�^zT��g�6�7��M����H!%T�J�#�3�����Ņ���
�S�Y�m
�Ӄ��$�<�n�T��4�4��Xq���)&́+>J�xf/�0SC��(R��秇����!�jۮB�՛V����_Ū����*8�#81FS~u�u$��QC85I"K�)7��Յ�E�#dJ�=Bސ.^�
Ar�	]�HW�0䞳��x��>�ѶrE���1u�3J�#�T�!����Z-�|�Aڸ��\�fZ�h�g��jy/��@V����Cd����&
��W�uz��
�c�	�}zV�)�����x� ����'�_h}((�T쓴[C�-����D��M/?�o��M��/����1��} ��%]������F׳##��t�U�qܧ=�GЙus�ܖV?���VOi~��f����?y=#]Qm�[P37��i�C(�+.o]�d&
~��S���_�y�ޤV���LU��#�b�R3�]�^�Dz4�1y9�	/�ʼ*�W$b!���bp�� 9�!}PK�)[:����?պ��^�/&C�x������;|K0(�Z�*t�O�tY�.�d�`���gf��(�ɸ��,�X�_����|3�2Ff�������O����� �k�B��+��3��N����ܦ����^����ƞ{ �.d����l"�/,� jX�`������J'<�9���D1�89���Ę��U�Dy0}l�	�&��(0>耞ș�F��K�<��]��$�����F��g&tz�ꐧ>�h�b�V��)�8K�=ޠh䞦��/=�	���ڢ��̻�k�@�AF�+�Ř��+�6s�K�(:�9���{R�kʚ�y7_bda&u-�g���)g��3W٤����V|�$�����+_rq+#���%�eP�q����xU���=w�b��u�F��2������q���z��ƃ�L�v�>��h�f�@)����f|�U]��9ʿ0��X5p�Q-p�Lr�"��}8V�y�MY�������U�>K��[�?v�1�4 ��CG]`B
��T���'@�Dd�m�+h����}5����\��
R��y�KE�~B��lz���.f�_�� �2��i�+��24ѱ:��@���>�8�� N����]�s�{LF�RU��T �M��8���7�;(�����ʃo��+%��"�"6Ձ0ed@�Y�����c��Ro��g� ��-nո�~��U�|���
Ph$tc ��^����}��"����~�m4z�3�I8%ϼ���I�k�'�c�̐�le�[8�s���.p�7x�)����-�1]��`���;v?��w�QcW�����a&;҇5.���#A��!�K<��\e���w�=:+$Ȋ�QП�D��t����E�s�����%L�4�/��%����Ы�OƖr0�s����`B�sY�B��r�x�L����y������Bq�m(�DȮWR�n� ���Q?�ݹrƒS.\m�4:xs��#����b�FEۯ�WY3J�l����{#�_P����ێʂ�fI�+��`a<�}~�R�f���Eۦ�V�X&Ň��xOn��u(��@�A0b�Eh�b�gp��ۣ��S\xU���8��f�.���G�~��xl!9Pi˂�J��xu��3{���D�? �@�������U;ۗ��g��k*���^��H<�(�� �H�<u&���]g��9tR{B��Gx�@	^h�ӈ�[����K����4P@�k��r1� t1kB��u��'�]Qc;��T��t�%?�H{�s��0eA��n���b�!��c�^F��Mk(�P�r��;f�3�����4�V�TϬҦK����8T���� D���wfςb��K	�㈬qsaaT��-���b�
�]	;Y)硈`�b��m�3�y������s�p`�ɬ2ޠ�0>�����kZ�n�	o��A#p���St����%p�g+�J�3�}7�/WPV]U��e���gOW�����ZW�:FX`;��44�m{�I\�������<�R�%?.��>��f�4�*@������:�����/��6�aRo���0����������q�
���&E:�<�!e�0r'2���t=���$RWإ��*�,2r�,b�ՓW��.�D��e�c��]qg
-ݶ�)^�9���k���I���s�D�ٞ���J��/<n����|��5oO��i�d�4:�R�-dq����?�3����Drz6�9�sc��3Ƥ��~P�ڦ�ze@��<��g���s �=��igj��M��*D�L���_�s��s$�O���B;�d�C�1@�{(��$$�iE���֣%����ܿ
m����<v�
	�x����	��ާ��3�3����ٝ�bO���My��dY��J�AΡ!�*9�A7�+�m-X�)�\���gz]0�OC9A�E|}�<�א����&��!���¢�}s��#�*:��w�-+���;a����o�~��F�%����/�ׄ��1���sH�f}�;�� 5è��Ne�g���1����0:|~�� m\����0�؅
9͕+�{q���� �K/+��;������:%�%r����(`V	�0����Q��5��_x]Y��>�'���<��d�j(�g�����d�J��/�a

�gk׾�E�w,@@Z����m��ȝ�~h�8��֬.��*e�H��c4|�+h�z�*��gi�Q����ǋ�+�Ђ!���|�� yC���D>A4a���G�}����s�(�H.>ڎ14 e��e�9�^x2%�o�v�Q%�(�K�
����i��	H0KI��%��)��?\��E.�c��&Lu��Z�"��`D5�!%��8�>_ߋh����[�V�����B���#�x_�m��VV�AgE�K�w�D!s%�δ`���D�-�޻]�h4�`�8 �t[��k�%ݒE:v�|��q_Q�_�X�������w�(V�G�!���!�l��Cf�(�y����S�s1_��Ad6�kY3
��g�K�+� �AԠ�`���>;.Ǵ���!�:��_������H3*��N����p}y���+����x4hI�g�q��j⽑��I�SsPo���հ��LC�t�Ԁ!�+6����{�^��P9u�:���P����%�RWƎ 3��o�/ڳ�	�p �8%��*��h+R�+0��ɡ��[�3!�cH���Vc��6h�МD�{�����p�+W�*���q{$aHi^�������ҷ�`����(�t������Ųk�|�<�ە�3�G|�GnF��"�N��89UА�ࣱ�چ`U��ľ���Q!Ām���Y��ia�<y��l�Pt�dB;�c�<\8��q��U��%g�	3�!~��H=	ӝ'v�@���&����s��H|������-��E }']Rz����3�L�_���M�ԇ����c��J�`��i~Ҭ>��!� ���1�,@���^S�ǋ�ϖ����ph��5E�=^X�0��H�"}��w���raM��������&��	�ۓ��D�"��Y&���1�n����4"�n�NE��w=���JߙV?h(���<�I�A=�āU���6��H�2;1Z�k!v��6�3d$�f���V�ʟyC�׍l�Io9]7j���Y�*�<׻T�2Q���c0�a�t�EaG��k��P����'N�pS�����8�hv"sk���_Z�V��aa�'f@v��$���7�&!���+��~i0Q��(2ΖD��&���jK�}�܊�͓o5�s�
Amn��nE�<bv���~k���A�8a�#�j.���ʌZ���_����Iqި�\�6c'�r�}NѨ��]�t���S!.��D�s��hp��f��ֹ�����y�2 �h35�t����K'�=�M�c�J��K|��y��ͷed�	v˂c8"B�?��Ƙ��a	����1�H��X�H�󐆓� �'{ń��-<f؜� �l4�wGgφ�}O}L�C��Z��_�9�ڃn��.�{'��ډ�� ��3�g���)^n�qz��-Y��T=1O9J̽A��-��:9E�Ȟ�i �*����pU�"�竿���
���y[���l���齗5�jr�&��	����	+�-DXf�h���"aV��[Ke}�["g�� �A�=���� r�
?��y�d=+ZD�6�Z�/g���&`T.�1P�l_��ai�_�my��TA����'?h/���0Rp^`.t�����k�f�w�ߛ�h�i��	���}�X� ���1�DS].fKє1�g��T�l��1��&ro���&j���	`Ȍ����}c��Ĩ��\I'��!\p����������V4��F#c��u�)�J��l��e�A�	�1ܻ�a�[�}�tߗ�<|\�D�ظ��j�*��.�mV���Y��v�=�O�/A,�eق1�U��G�$�'o�Zo �WWx��͠�1�V�i?̘Tk����K�2�r|�W�N2�Xo��:46G9o�߲��#tŖ�b+�q�P�)�[MUŦ�S��H��}t��H�d��-�'g#��5���_ $ !�5;��TXW̟�����(i*�p.��7�/]��%2�X�"na����o]�Y;��hyx�o�����q�:����@�k�:�]a����o��V� 1I�8���ʼ��� u�DP���J"�	 m;�Y��ԩ6���l�r��x2G Ǿ˂��3ZV�>��^����(o����`sڬ@5Ԗ��$�%��a"��C�I�}(D��#�������A.�����A
���sG8���Ӱ���K��UO���<���ȗ#�=C���MX��y������9@����b��&# �9�Yw����%��>4���ң��I��'�ed���X�#��!�sL|!�����+!�6�)v_����\A�Tv:��y���#F�g�0�Qffe�m�y/�G1J(�F&�S�v��S�����xn�;? �6�D�]ׄD�