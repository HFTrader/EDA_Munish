XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U}��יI��H�5K��>2Ծ+*3���I:M�V��a�M2������>ܺ���'��%ĳd~��o��	ɐkw�Y���*~��h�����" &���
��Un�����9�ɏY�$�J�������|�m�	,@K/�S��K�-��י(R ���4���w�i;O�aې҆�:�Qa��CN=0����ɔ��<Wǝṁ]��l(�d�LV��diw����w2<�����7��L��v��j�kM؈k��/~��ώZ��ww��%�D�S�0
�7�0���q����~�{0�-vK������8�����NLd����<e`F�'PzV��rY�~�H3a����P2�U˾�,!1��C�P�V���9��?�誧�b�/�.�a�x�����{�`�:3��m��)�a�Q�4���9�B��%���*?�C�>D7�S��N���D����g$�8[��E�m�&!7�4O�)]���c'k@���凹��;=�c'M5y�2d�t�U���ڲ�=�S9���#ŊK�"{|`[ǽ�$<���W�*�+6�p�ܟ�;�x[�� qD�c)������#R���z�{1�f�x��X����0!���7[x�D�A)���5f�'�4aۤ��o�5d��I�d������%ny��������H�����>!��f#(`�8>��Ϛ}[���+��LUH��X�6Mnxޔ
��W���n�(���oly�ls\�F���b�����R�PS����<J��XlxVHYEB    5e2b    1530�7��2+^� ���_�Ezϋ�]Tp�^��ȷ=J����ϳH��o8��<�Ut��Ё��R:@��}o�-��ͬ���/9S�pL*�i�"����A
�6b$�eZ�jz%Z���R�LU��X�my����������,��R����R!`��x��U��wƸ�5����jO|��AT�P�rj�c�^�[צc�c��zz�}t��,�ړ�4:���?��da��@^�{_�kVB[o�S���� W���儣a�;�b�tbb�f�'dF��x�I"c��{�2]�Z:���swW�S���0�88rҊ�@k�{�oJq�-I�O!��sq������D�*A8"@4�}Y�P�'��)l�*^����a�o��}Үov�ͺ��ϲ��_בk�!��a��6��"��9����m�7
J��2����C�	u�G.i8� �j0�|��2��Z�(�����=X�)d*l�WJ�u/F��p[����̮�K��ͯZ���4E�,�
/�_�-��Ặf��3�`h),U@���o�����[ES�>ŀ���J�\Df�i4 �����ϸ���^s)�k��HK1�t����V�Vl��i��w�6���_�l���8w��xU=�_���&-��D�2��{���	zD�ƊK�"���8� ���h{���>��vד`��3XB��\�"���Ҫ�o�(�a8Ӂ��"�|�+�霶�i�OXˇ�r���к����l�j#���7����r4�O��������y} [���$'��>#|O�4��[�S1��K�3hR8�b���dѣ�:�x�~ٿ�ON���K9�/��1L��a3���pbZN�	�����e��KO�w��8H�g�y�"ʟ-�hwA^��@���L��w���%��I������ޫ��&��Z�_pp|��?԰�Gw"��!Kj����~V�L�H>�w �ʰ�E*ղeЩ�%1#dOL�'L(���(��m���u��=��+v�כ��c�mw]}��?L{$#3��@�C���m�|���p�>TJ�9�P�6mճi#G=KQz�&L}y�s�Jחi��q���4�����pnzE��^V2�lu�r�H!V��[��y�Y^�0d�Tz�&i"�2Vȓ6>t�|��b��X��7.��dJ�%�&Ɩ���`yWig)��ֶ��}�7kt����+�`���Q�K���>�w�8i�g�:u��&����y�Ю��� �,�Ϻ)��jWO��^��Ӏ4Q4�"�B�euS��a��&w�O7�e(��~����@3����9jz�ݗiЁ�;�m�Z�À��h�\\� TO�1���,�U�&���.�q%�W�=6-�("�@)J W����0c�J;����g����[�]vB���S�o�k��$I��h-�y�U�$Tc���O~Ĳ�6=�'�9�I���'Z��XH^�W�6�6h߆JoP ����e���{���>�u-�A�AK����!߹;	�#O`� ��iP��'&�	3�4�Jn�(G�R/j�)�vxU����`[J����u��o���%��;�/�X�(�mJ'��RP�C9�}m�����W�PH1�Cpa�p��|��E"�S?yv�%������v��Z��F!՘��wJ�2����c_Ƙ���e��/a��|�C	]��wGjk9�Ùi���w�y����
`{Le3��]h,�b,��|K���Mɕ'cVnHX�H׬��uڰpt�B��wka���]1��Y?ޠ�l�JJa��u��PcX����+c읧�w����o�L��Q�.�[ζv��j��|�u���ɋ���q:��z}�(z���d���������㘇v�jGY�6W� >e2;%#���%�g\��䥝�-�����#��J�ՙ���?��j.�mIo}/�ib�;F��D��e���cn>yx�*����q�>��z:�˘�z-!ĎApxr�& v#f�4�M����7E ��?�]��|��{Y��0$>��1����N���r�w���X0L�(�����$��9#�� ո�+�)���t-w�bI��l��室��[��-z�KJ�Z!G�� 䙭MBީGa�&ċ��DJ�W?"��s�(^s�etG2��\&{F�kI&
s���e��P���a�Gl��y}CoEѻ���zww��TO��&����/�V瘱�B��!O���8��L�.R��+C� ǥ��䉆�,����ʅ��2g0�i�Y�c����/. Y�S��į�ѩ�ڭU��/���sQ�k�q��J�O7 �/�3n-�������X�+~�8О�~F~�!�n�u�Éz�����Ɓ�U���H.�F��(��^b��@?N9�̀�����������~�Q��9T��[?w��<́�V��I��@�)0x��9����^�}�l�Vt�c�d��Ho���έ�̄i�&�����t����/���4M�uE��l���a-2�������8/�;�ȼd���H��Lm�}�/%2� ؈�
�DXm����Y��}�q��a�om�+�99�X��U�Qy�M+��,����|�E���/z��^6D�p{76P9TU��( �Χ ��q�����n���/Β�h+F+�\��K����f�=�������=i�-M������T�"�X��U���W�T�Ƚ:��"�������h�)準);l=���9��i}u3F��GY�>/�P(t9w�!'���wjE��際B��W�p����~��q7�!C�|&0�䖆 rg�iJʼ��ʝ|�O�^�؁���q����Zuj��F�. (�\�� �F���iZ������f��^�Wj��9����L5 �J�N�Ob)�W�'�"U9E����=~'ܷV��NE8�T���;�~o��̅��e2}�_�ggN�$���|MGV3�Fsۥ���;���LL�qP@��}���U! Tiyݎ������3�^��2�O�����Huyֵ��ܠA�1�jG�,a��K/ӂ'ᔄA�ʫ��=K. ���	����E��1�|�p �J�k2P]1ׄ�:1���S7U���'b%���������[�R�ך`���0��@������.�ͬɻ��IJ�Ȳ��ƙVZ2�uf |��D�Pj�̨�p��4���[��+u���f�{�tp�p1M�G�C��̇	E/���#1 �6���H��SO��5�-rÞq�v0Q۫$��,��1�����SD&�^׷�,0�)��d��8*Yj�Y��)4Dl�=�μ� BB��@�m�Z*�NL�#�}��g	^Pm�E���f@Ͼ��1�<e)�ti�]7x�C�CV�L�(y�=J��Yl�ׇ;C���(/s!l
޳���·��⋀U�e?g#��X�EI�%m,�͂K{��&]�%�+J"�V	<�\�27�'���T1�v���=P��ݑ"z�ّY�ѡ����S������ɇ�r�Bf<%� ]ɜ��%���&0�{E��֛!�{�X�݄�rV��2jޙQ6�>K>Z��kC#���D  7��AA�+o���.E��h#�����_�Q͜{��� *���Ɵpw�|[tA�fk�z����P5�
��ZZJ���,����s��|zt���q�,{�?��u[��8�-��矨l�gO�DP���~�|\,�cZ�"��G�n�dƕ�a�6�YΪ���c���>�&�WE��j�rcSK�wH-���R�3�.���x4(c��Ц�w'	����yr�v�bB�{`jIB�?'�L*_�-=xT$F�Fz�Er���@�A2'�U*���=2θ�|}��Z�ן��}u_M����eV���O��1ݫW�Ɨ���K₌m[	Ȁ|�r������X��ߪppT�;U�����Cev��2��]Z6� �`��x�E��R��������a�φO���nTC�-��~1/F��`ɘ)�ޱ5��zS��D�%�i1�ǔ�m/�6��Q��:v������q!j$0�/���-��=[:�+�NX=<�hc�����sV�H�A���D��XK]f��!�^����3��m�ܸz��̤{���m�$���	[<PJ�E�INlf������b�Mo��s�*��ib�x�Q��W��ƊR����
,K�7:YaW�����:�J�Hw��ʈ�^�2ȸ��>��2��dv-��%����'�)�2�pYt��8>�	bM�15ń��Y$B��h0<]˯�{�B�m�Byr�
���r��6X��eN���b�$Ё��XW���.�:�$[�5WTP�(+EĢ�\9Q��h� H����oK~'�mb��U��IYCC��PW��� �C���F��Xޢ���#���'jˬhi����{�2۵)\� ˣ����7u��+ܻUE�-��EN�s;
�+�@��åz�H�6�^JU��3Ջ*b��~X�H���	d��E��	�=ƹ��uE����J�x�aS�*@=��4�7���^f�@(.�sx�v7Y$�QPZfԒy_�����9(�uX�a�L?�@����t!}�_d4��.H���F}�O]cu�#�@�?p_�%	cE�<��˚�+"��΄���G��\Aggz4r�+������GuI7�0>�������*b)TȁF*'�X2���=d|���<����J���&E��ك+ �Kf�U`}���L�i�wBAd�OɸRt�11DR2��H��s��?���0�l���,0�#I�h��t��RM_
;�Q4ip]TZ:xn�_mt�\�L�ѧ��r��3���U>M����T�Vd�Y�W�J���d	���qm~M�B�z�dZ�uR+q�)��<XM%�߱���}���x;>L�Xi4���S�[���S��x� �6���4�vZM�ʛCRυ�F��@��F���� ��{)n���-xOY���+��=I-��^�A�*܎Nݱ�֮�QGڜ���1����Ҳ�g94A��љ�A��\���e�M��e2��FiJx�TKM0�v�U����R\�������j��15��.�؆����>��P��R.��G�!��}o�~pq�O��^��N������xVkF���3�_�1?]k�W{6���>�����Y�͕(�|Lh*���I+�|�znP��C*qZ[��@�ڱEu��!6�'��sPR��q^Z�e#�g(ct��ʶ�:�����Q�zX��;�h�t��Ӥ��f�Դ.�z�_#6q��\NȌ�4ֵޣ�p��<E��׭3�S��*�y�y