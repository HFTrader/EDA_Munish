XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ҍȣ.�Br�8�ܩc8�Bj*�(vyT�G[������K�>�C7�����׼^����'Φ�.s�=%R�����{(IE���ࣿ�]~ժ-@��^P$ƽ��zd;0?F҅ᜢoO(�1L���%��6����B��|�
Ub�!$N��:�i���K���؋���̜WY��V6�|���sn��/ Q�	�n���惠lؿ.$�򣩜��� �D�4)�2�q����������'���$`��/�R49��P��OC;T+f�b+���rЍ���
e��/��7�1��[���g/�-�Vc��/�c��8��_���	G"��nR`�A��VKi¹u��D�l�+pL]W?��/����BlZt��f{U�Kq���ݷ�IF(�9O�����ɚ������$Y������Sg5V��ա��%I%���^�FK�>�Kbd
�s#�����Ͱ�s~	�?�lj3j��Uv��{���)c��|rlha	N婨[Pe�س뗽�Cl� ��fv��J����3-�<ԓ$Ρh�UC�q&Vr�UN���r#�W��e�[,���jP�H�f3�3��i���W6O�F|񵼌q)��^*m�5�Ϳ}˖�].M^ ��������j������o�@�/L9���ź�+pjl߻�/1�6
�+{HJ��\B1L��[8�U9 H��Z�G�&�GeL~ ��.��zB��*�T���1_#В󿾜������2XlxVHYEB    66ed    1670A��c*z�F��w�%���x�Ӆ�7��7U0���B���8M�b5�K���,�7������H�`��ٳuuW�9�5�ѓr�#_�ھ�rr5Ȱ�a��Ǉ�����~M�[���ʨ0���g�Ȱ��7��G^�{5��E!s����j�8 �:FD����]�C�}��e?�v�j!	��¼�]�rJ�f�v�Adl�����9ȶ�dM�h՟Y	� �s4v�?�FX�;�7�I�c|>1�D��}M^�.c��m�e,?ۭ@�g������v{b}������ۿ��WXIe4��.����I��/�	��������Ӝ��C���F��#N,��G�%	���7�,���{m�.����������̣�t�wr��r�M?���b23�2����'ac�!�=\&�,�Dw�ݴ��-�"?��>�#-�3W}��7��a���ҿ���|�3���$��p}+���z,I��f�r����m�~O
M{��:o����[H��xX`[��7F/�[Y<�ݺ~~\�� �˿r)���@�3�#遢A$�������x���h����"ئ	��cr�~Ɵ��\�6B��jN���]�"���)�y���q�jq�ڢ��l� t��y����h&����[�� @7&ZCS��������o��yO��������\�m?�Y���ee���������Ʒ���<��MV?�7��"�#3!��sOcu����y�WnuK,�u߯��IS@PܒgF_N��.�dr�h��{#�ݾ3�*��E璙jZv8�c�F�Bz=�k��5*3��w��05O[*OK����I���6�;�꾑W��9IF���I'?�	�1"�� }��u��1���c�]��Dg5��-y~6��k�H!	�lڈ��{v��͏ ̟J�L�GK+�N��玝b�qd8��-#�����I�4�yJ��r�����vl�ߎ����ȑ�(��]??�5%]@����4�n���K/��d�╎\^, ū��&'"`�����V��U���C��oc��z��i��P�&E��]
���5�l7��ΞoaA��K� n��-�؅�̀ק;n}o������c0;��M0�@�%&��Q�;bWW�[̢"aݓ�݁%~� a�p3�eg]���#��֧j�Z ��=���y�nd�V+����%A,(f�_��y��)�Di�w�T�#�בU(ٴ���%�+�!mN	�jv۷f��kG#��䬋��-�"N�����RZ�ϩY;� j�2��T��3��F�|��:X�3�Ch�ƹ���V$��"T0*k��x���x�[�8)1��� �=�H�g��V�\���`�[ N�r�_��乹��V	la�QwJEn�q^����U.}rL�Bܒ�x�mp$~�O7d���Ce<�ݬ�o��!�]4*+�f�a�Ӛ���V٬�_DK�a�c�J8`�aN��eCN\���5�s߁��	�i��~>��,�\]D����t;՝ε�E�ɏ�`��g×;�u�X���K��g[
Ϥ ���M���2{L��p��$�Qx ZQJ?����>|n^���ö�r��������ա�������y8
�
�>�f*�C"U(.��Q��}��]�4�÷��<k��t�H����ta�1�<���g_�S|e����hƉ�1%�l���
��2����-�V7s`��zo$��y7i궱y/�|wT�ă�x7�ہ�S�-�A����OW)��Ƽ�g+��-�� ��x����T�+��rG�=Wn.kN��ӓ���~�BA��8���	I��T�Ȏ���RH�>��	r�/'�.���~0�w�;#�g]�.2���ysW���79��(�;�52] �b�7CY�cՉ�T��jBeX:ϧ�&�TE")&D}g7�қx�0XC�;��F��m�А�Zq�ڍ��>��辬�6��c��U�͋��S6����6�L�$�s!!V9�(��=������B��ؔ7e���^F�A�˽;�7����$��#Mߨ��9��-r��ZB�"��UG�u��M"ބ�~��� y�韷�y0S��B;Y�"�"2����eRm�����Q��u1� +���+�8hx''�s�����S'$L��EcE)��j�`�����xlr|��y6�巓�t*�OXԽ�0�������K���R�]YPv2"�t#��*$�T��I_�7"�sa�i2�m��B�NL�;�����&	��:�w�f����rjoX;�'IMU�bͥmI����2H,��������$��ɾԨ�Ę��4���5qP�7���ڧ�k��� �Bk]��So��T[�&�췳v�º�jd��p���nA���Ȃ�����1a�X�A'Z�8jJ1ZH�ܹ�?��
��K�<�/�����'�ϐJ�����+M�4��c��͹4<��ڎ�?5t�e {m:+��ɬV��:�0La�a��%(Uh�b��)����1#7@+; O����!y5~e���H�/?�A�=�`5���Sll6χh8�~��UGo���QET#��	+ �t�)-e�ŗ����KA�X��"��	vV�	����'Y����vĕsP��������I�Eտ!�� ���P���IQ��إ���t�vG *Q��K�K �w9��L�Nܜ��^]r�N0�~>�'��G�Rn5��fE?Ȝ{!%��F���ԁ+>���7p`Ơ��o1���a�}�n��>�=H��ť9�uؔ���֯�L���*[����zrM.�Y��9X�u?�ĔJemH䚸��x��Q�b���W�����j:L-@�X9�ڽ��v��H�����	�.��Թ�&���;!M�|���R���$�EV��^��<A���p7fUM�q�������T�fbt�.bF�(Oy�����7_է�\���Jh	<�S(0��o%Wl�c�c��2a�ԷW�$��2��d��®���#����2��̋�L�������hs���K�.��&�߽Ҥr�^�P#e^`��S,�%�A��{uIO?ąY=����H`x�=1���g�a����!^p��Ad�A~�����P2��,��=���I���~o�����^�������t�v����?F{!�"(��v (ǌ�@�G���-�4N��Tۄ�U�ڻ؁�Wd����1;
� FDL>�}��TXĪ����M�7�hd�!S8�]	k��=<�)���$-	LpV}�L����D�$놊�K�Gֲ�����ݬ�����=��z�m��,�r���5�R,[�[p����j�u؄C^��K�!���Q���@����U&Y��5Ⱦs�rUŃʻ��A�'1��D]IjG�
n\(�N�Y1�x��d
#��܍^ztֆ��j:�l��xU�XR�v���6�@�7ŠN�NF��A�'�د�Mz����yhq�<�UCrO�g�P�Jy/��|E&Q��t �=�o��e�(sh�6� C�QA�X��
'N�5A.B�� ��6^k���R�;�(�N�j��Q������V(Zx�N�X��{)�M�n�~�3hN��S�Um�i�=�M%�oI�+�nr����#z��\=��lauT�ר^��T�t>@�����	������f�`m�	�TY��&�����C�)�!�t������iVK����:2��j��m�����j�O���V�);H"1s��/�Iko܄Q�@�	��)��'�O�����}�*������?G_F�뀻'q�@�/4�Y����*G�
�W�&y�c�xz�.i³������3�^��FjmF,Z�8�v��� AV����'j�)�}P�$�s����� 3��A\L��F|{[���F�T�m��!�J#L�Δ{шy(��XB�J"T��F�`��wr�];�j�O�i��yN�az��<~_T��4~v��#F\N�ٛ+=P��%55���K���k���Kl!�*�#6��V��e-��i�����NQ/\%����i>�bg{B�s����X9��Xڲ�I��_��B)vϴsD � ��`�ߒU�"��1�0sڨݫ3�si&����!4��9�ܙp{��H@h����=�/�X���n�;�/|߿��=fEg��yV߿!)���J�w#o�Z!#JX;#;���Q�<��Ky�A7����X-*B�?'��`nu�o���*.�%ɤ���|#��y�g�s-���@/�sRO��q�*_~�� O��>�	ʧ*���U��(ˢ���; Y�ET���k������V�F�Df`��W�x��T=
4t�A�kq�I�$Q��L�Ie��&�6;WBTM���El.��������נ����&�>z�1Wv��Ck�K��,� `<�=+`�-�hK?C-$;w)��p�8<���*�@lc��W@�����\�r��!H~8�Ë~��ɹ��--���_($G���):�8�v#�(�BUh�R����vL�Arj㈝@$׼�$Gm��%Z��b��q���p��[������o��(gȄ/Q�$
��c�pF���*�������Ζ��6:��H{�V��w��nNd��T6��nЛ��a��q,F;yߨ������N�.���������-�Z�U	0B7Dx�FG���l��)&dx�2� $�.�"fD��-c��-�b���)����؝�z���>��V��خ���U�������~C� Ov�0�b���yO��y,~��`�XVX8/TN:ݚ�`,�]mmt�̺����5vD�j-��fM ��n�O�}a��P���(���#hkx��Za� t�J�ǌא�/xM�y�>�5�
8(���"V�ߩ}+���QjFu��ⶼ�|�;����u��C�I9㐴�`���י���^M�HNg����{oI �+6<�m ��xsz�mĥV��ۭ��pC*2I�ˬ��5����&��x��{0�A�YBR�-t�b�>>
a��J��[r��e��,�!B���;��2�p�K�&�S!��A�����>���W|c�� �@��s�E����~6�����[2�4���22����#�"l$����>t}���&�slv�����U� (mBjO������*��s3W�~�~�65�(�Mg��6S���k����j��ph�/@�N�Yh<�� P���e=�Ќ�6��q���O�*n_8!�a���Km���#���P�wq�Y�=;���Q���E�h�c >P_���z7�槹a���:B�������|��pn����	�y�qI���Eă��w���������:�+�p~@(9��7�E�+ߎ�	�y���He���_��O�Q<Ͱy�g�+엀1�{c.$�o���<1��i�Z��7��
�������8U6�`�3m��zI�Q6g^3>��zT+�"��al��aW]�f�d��[.���q��Md@��%:�(c2���3����~�0tB����>t"}ԍg�Y��C=��]��s����'_;z0�m��f����x�f�H��"�A�yk���#���A���L̃��I��\�l��T�����~ׂ��໨��ȋՐ���Bm,}��1��\�<t1d5�s����&�d������x