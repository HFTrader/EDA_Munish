XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���¡�␲NL�?,�J�����s}Yܼ���s����9�Ln}nǄ�7�?,7C,XW���ll0���L�!@�@G�6��}���-�D��,"�f�#-xKѺ��W�|���� ���75�+}�$�y�X���)��&��E��J��� �*a!	�n���"ϮKU�g�'%/c+Ӝ��jJ�D�r�Y�7����q>��M⾌u	p�s��͠�h�!���,s}�	Q���R
��ۣ�')]*]�<�i~ָ���J��L�%@���5�	��ocj�aùC�%h���\I�X{�n_�I���bP&��_lk�� �,eS�g�E��6�H��ڮT��B	��n%w�%?9B������.�p���ߪ�w�~��H�_�堀S4|�oyӺD�F�d����� H2ԙ6q�D���ߙ�m5QSE}k�ϕ��[���Hy`�����i4*U����+=�-�}a��3����Y�Y1-Ӷ�u`D,�����(O�F�؜�c�B$�ͷ���Y��hњmf|TpR{��/���戥%��g	����LH"Y����`Ȋ�.�ͼ����7�%��K2�0	K�5)o-�^�hz�:�a�'q���J'Lnې��^/WW'�/����tWs�K�]���~�y1Ri�m�	E�h��7@j~��(�X�G�q�kH�  ::�i����f]VvmgiR�RI��CdbG�p�q�/�N�uG��r���`'�]~Z��K�^D$}����V`LQ.$�&��QSu����Y�;����``XlxVHYEB    25b1     b60b)�Ďwlr\!�����`�JV���\���r��\�����t+š-�YI뫁#|>6�,��HX,=�5��T��o�PC�	����a�]�l�t���f�&�es�-$x\T��Z�Ҋ�0N���T�U�PB�VrP���X<����~�T��Մ���Ϗ�����Cx=ڔ�
�${D���������
h��w��;�xS�#3�~�@��� � xҊ�9r�eY���n�ų6��z�4_����cAȦv3pO���l���(��w��Yt�<�WP�l�Џ�|۾[�N���s7)�.�=C����ƧMJ|Ś��Bʍ�K\����vǃ�H�[���&��&�6�>��N2N.�%��w�����p�@ �<ò�\�K����p�սZ�=��Gt�E�`SX2�h+	O�*v�Y�@�Qt��gZ��g^���x�]���-Y���%O�~%�Ɲa1���	�/.1Y��Lś��k�@�;mSn%��'O֋~:��e�$�hgw4��Yc���ӍJ���~&|4��9� &E2��}C rR����K�ƪ5;�;��񡮺�$Cۚ���_���Q!��?n,��/LH�Zi��C,#%Q�A��k���M ����.7 ��[���b�L�/~A~���Z��������>�c�c�F�����Y
�7�5.�&����T��E--뼢����j=��p����9lQP��F;��-G@��ƻ�Q�S���Ĵ^7=X[b*��?�c�(ν0'�L��HXf���(w�:Đ
9D���#X��7~T�D�B��8hz�+�=�B��a'��0a&��B�qj.w>�EɅT֣=�C�Q|���=�	��	���A���`sFd\�}�R�wTi�|@^tJ�&5®����6������K𨷒�?[�%�3�|�`?7J��Xm�2�@-	�W�š_�D$�A�{ǐ&F* �^����~��_X&��>G[=��	���ďO����V~��|d�;��s��n�*��e�л�:�g���S����W�2@����3���@�ɟ��[�L��U��+2���<��k���Il(�����l�
g�^�?Ø�tK����纕���4�ǆ�oA#U��s�5�_΀K���/����8K�������]k��,�/=�{�	��!G�� ������S�ȟ^C���$1�3�}��	v�r-tң�
w2�\�mAp�B$:�@�"�r�[Ŋ��;�@�mv�g�_�1�b��`���t2`���t�}��#��f��ūKt~�c�=�Zۇ� 1o���/�8R����=fS�}�����Π"��}Vy-=���kh��Z�L+T��0�n��<��(�fY��:�o#~'��~�%<�����,��=�W�	Ӝ�>O���wI��C��uJ����\���"J=N����qj��yT=�w�q �Z���������1_�gWX��}����HK��ݨ7��k*�q�m��1��ŸHJ�8�V���匆S�1�3}<��,'RƇ�p��#���6OK8�"�\��
@v�6��#o��)ٶP[��C�E�h��܀��zm(7ÝN���^D�E2Ūt�Z�?SN�����T�mO�9Ϻ�|�Lđ���Ѩ9��N�N�������E��û��{L�ͤ���k�s�9��2��Ę2]".�,�I-�l<ooj_YM�P-�>���i	�J�߂��B(��LZ�n.��s!��0�@��%��R���~H�J�_r�{m��0�&}yE�ϔ�ُ�/f��U�}�K!�4�e�'�su��y͐�������6r�l�za�-.���&0�κ�����E*T��lۚ���g�� y�p8hG;���X�w�ߦ��~6��l����p�W�N\--*�i7o�:�j9�WX��n����t]v�5y����4@��N�	�ɘu�|����V��v�=1�_�Ō�Հ�|� �Z{�e�J���߄�l;�Sl,��ܿ���^�{<Q�B���B����8�}��wmr������*T���쵲�Ԭ+�.&�;��3�{׈�dߠ�n�K�Y��VW�3�
k`�6OF�*��$�BY��˭�g~��.���_�~ݚ�	z���L���<+�D�5-T�U��Y32@H�����6g����
��h'*8��bQ'wS����*��1ƅy��|Sm���d��ה�m-߁����Y��Ѿw�=��!��@��� �G������k�Z�3_m�~�^�	�ڻ)P�1g�o���ps�-�90a��	�؟ċ�E��G��#z�h|-j=t��8C�֘K	�ˠ����dڄAh 4��b�7�>����~ۮw0��Q�bC(���~@*"P*OCcM-�,�v�@{���H�-(5�iQ<Э�Q�:e|�/�XKq	��{)�	} ��$��ux�Hiz��t~->�PP���ȣ�IV��������X�l];�&��2"w��e�@~ҿ�DǶvD��>N�D�7�ӋU!<�y���Y�*fY����ӥ^b���a<a\`�����R�x�b�9dZ�X����#`,�^�֘�� Ν<O>3O�ӷ
*p${�(���(������>����'iI����A��7�����ϒ�� �ޔ�!�D�Ɂ�5[:wU�"8w(&'Q{->��AuO�Z���?��r���O��ܼ���̟ֆ"&<��u�~�"�wN��BiiC���XԲH�V`� LD;�R8���5�t��x6jK����{�冸d�<?N�`Z"P��ڕ&�50{��w�&*���k|m�-�ć5�\��Z$7|")g:h�>§.���Mo�1�L���{>�a)��