XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��y��N�����V"+��A+ר� RkRݚ�W|�L�9r��}��*��PQ*J�L�r��"SR��+�>�Y��g�3X�K��5B!L��!�^�����/�6��ǅ���褚�#8�M�g (+�<%*&����F���L�ԺII��4�GAH����l�ޯ��f���������9 �t��9��B�#�?����5+�r0�?��,��0u�)�A=����2�� [p�};��!�&M�T��"4�ϪI͎��:�i=ީw<��
�\��W�$��<F��J���`hp(cR��>5�Ӫ�Y����ᵄǻ�D�`'���s����;I��QI}���Kq�P�O�z����sy��ʠ(K6^�ZS�;!��-z���V84"���j"Ȯ-��c6ޯp5���B(���0����	��(�*5�����z�j8�L���g�2�b�����i֠��g`�9�v�g���(W8;Z�hD�H�^-�>�g�y�����C���M���/gD���O��/y!q:	�ٌ���"�*u(&}���9°2P�(䗨:�6kh��*h"�L�?�Z��XG#�sĜ!e����/���1�n��B"ɸ���`\EL�c1d��E�l)0�@R.�"��\-�#���E�����Q��Zh1&�X��bH�2��>�c�.�v\:<�џ�eJ��7�ǌ�ey�/AKQ|�s�:դ��50q��g�B�hteӓ�*�L�XlxVHYEB    1aef     950G����<�,��%Q��/SbıS!vs�SN�F��~� h`.�������j6�x}�b�N���
��f�� x�A#�7��/.�u���^���N_(i�YWk�Φ�\��,���^l�Z �]31����v2 �����;�����]��./���R�ٹ��9j���Zu��gA�^���-1"��@�P��wDҢ$;F�����*�h��U*$K�-�(Og�6\2
��b)�+\+�x�]WDr�rNR�&q|)#��
`.��`s���ۋ>�̿@�������G�eh����њ�r���4N�fK�fHT��a�e�g0�N}
|�䥣ÿJTBs��E��O1����^�G�N��-�w����O�1j $v�K�=�B�G)^��[���B�W�F����6$͆�&w'f�ic�h6�#�z�
~N��F��D�g���dB�#���w���
@��}=�1�P
?���� �����[d��F�SJ�:-R��31�<���"�;����܃��
 �y�@�/`��dSk�=�ubEK:"?�r(o�G�X:'��~T��3��
�H��f�<ͺm���V]H1eJ[
�at^�89���eS��J������.�z����*�����19��Sc�9�N�#�����-E���vJ��b��w�i�ZP(�o�@�f�{�ZE��A��@��$�2��P�0�aC����x����-�&.�.L�Y�.�SE��H�����'��ZuT��H�48"I�dG��멷kZ֪}U�����c\Ҡ�K.dq�UtE{%X����Ob��njL��gϩ*͞>��p��#@֞�^0�'0��K�4�.��T �,�� ��;#
���w��H��톡�y�7B� ��é����P�*�5��sV�D��,F�ά~�$��'����_9���,7�\�%�:�X~4Ý�g$�~��75������Fq�?��4?F�����H��e���^�04h��|�!Ghb
urW�-������S������f$0"��[�*��P�'�����H?�n��#Q����u� b���+��2���#!�`vl�?Pv�KS�2<}���L珠K��+R��\��sR;�`8$F���%�%t�/��[Cn�n�5��+�H�T�E���]/����m�iq�$C#�bu]�����Ŝ�q^t����6АdO1��Շ8�hR6T|�S��X�S|�KWal��URv��K@8�5ꯂL�������p����)t�C�!Jg[G��Z/�@� ՚�o�N�Ǵk�5�~�	�b&�O:1�w�PT_����7*��n>w���=P!P�HA%��0��Gܙ���:�-�U߱gc�i�	o��0��փ���e������{�H\N�s���EԹvA��/��xL��'c4Ms �+���챑ȡ38�VCy
�ڲ-�ΛH�c�5����zg��a��(H��YK{�(E�5 ��Az%�LȘ^�0.%�A3����H͗`}5!�)	�HfGW5w�y�C��\g����̬r��H�G(���E�����}��x�;������"��TJ�Q�E��-��v�A�Q�Q
�7ڡn;��4[�yF��lF��?�`vQP1�xy��/'�ւ��t΅�(v]q��a�k����X��q����T]�@�E�^V���S��p���B��@ъ0��F�x��S���y��A��Ve�n�+qa�P�����FΪϮ_15�N~�
E;8!�3��Ì���&*P�_퉦��1�K���H�<�W�� �M��Յ�,|�;F�c��P;�F}T����طYv��t�fR�Yt��b�g0�'8���g�&K�R�%��H9�_����z�&&b���I*��VnW�{5�>�����&p0$����K������9��������g%�k�?�,��x)m��9����[a��(��l�,���)yU\��T@�F+Z
����c���:�5��X�1�א���Fj�L�(A�c&��L�!1�O�N�-��Mp��߸%	���/
W��8��
ʒ�j:�ѯ�������)8v]X�%���'.��Nr^l��X�k�[7D�T�#�gP�[Gf0 ����6��&�Whj,��.7Tn$L��9�8�Mb;�xn20����I��E��yv�����:囈��J�$�_���BEh[:��H�q7��n�>��,��m�g֍H�/>�y����%2`��s�E�^�;X,y����Ji�r\���h��� c6��U�LP�HE�9��T�"���=	v�?��WAI8��s��mq��c��VhrvS�GLml6�9�>��ϷX��bVl��i5wYu��m,±vf�*�;O�L