XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/l;��RT�_c����ٽG7�����}e�?=�̻���D"j�h����KdW,ȵ'����z�n�)e�;3nt)C�y�[�D��L���rR�k\������+衸����Q�
Ï2L9\�Ùոa��e�7�V?�H0��T.�Y�L�$��D@���a)t������W��ޫ+��g��%_g���w�L��%�6�5<}����2����/����'/�+m5%�9J��y݋��[���v�d��b�;|=�>;T����xL��!�`����ɏ�O*��+�!�~
ћW���׏g�3����
�O?\�f�Y������?~������F�!��Z�/�Ni����#2�P��T���n�ў�*�*���>]���qa��F�`3]���3	���T$St�W#�f̮˜��(�ꝉ��q�p�(�*v<����]ְݜhc�er�X��z�M2��µ]�h>��B��D��������aG���KC)��O�b��A�$A�A�z���?�&��(Pe@�)�Aֱs�}���~��E���2�SCpx�ZɅF��K>{������YY���̝�8x\7�7�P=C��l�y[ |�}���l0χ��r���;�U���<�m�a��	���ڃ�$B���R����M�<3�N `%q'lW��d]��l|D6pv`HS�;��V�z�����-�6���Rأ@S(Lp�].nT�B��on�Ts�;g��) �h��*��24P��XlxVHYEB     f6d     6f0S�Sl�Ω,�V6����$��^Ӈ���ֱk8�[��MO,��n�9䓂����b��`��I��]qex���uLN��<�h�پ��7�r̸�[�@xv��ѢX�c4���M�9>|#lNؤrh �gbU�%w�
9��(��c�f+)�u����( <S�m{.0�"5k_��BkR����'L&���M(���۵���ۊV��1_�[}�\s��{�ab��mTHp�&0yn+�$�Z�N�)�Z��J��:)��A��e|A���M�8��BD���t��&�pm&�ޞ[`*&B���~̵x�k���e�=7��8aV��<�p�:=��Qt�̞L�x��b���i�Pk���̜ta~�2��7��;�Ӣ���Qː/��[�
k��3��V`�8Z8�c#'���\�I7%�=�gQ�& �ef$��F �y�+~n�@�62��0-6��]O�Y�Zi�R�Pn�آP�ԦI�:�]ů)d�޽�~)3�$�-����I�� �$�ߌ}����1�������T�rC��x��A"��j�_J�f�A��M���5}�*���\��љ�aB��fՀ�繜�z�\����K�=���g��r�~@�OJ��棍����^0� ���_����A�!��7`I�MS[C�!B�~�W��? ��|�]�Q˼�Tkg��=�!I+'��$9��?iW�����C�T�Sa=�wb�����2-�1�9Kw��n��¸�8��3kr��,�G�u�U? �炙������ی$�E�j���af(���+���� B�	��a�zd��Ug��w��#��U���R�~����D�1&��m?�Vy��[� M�.[�.c3�u3g�?O__F�R��uU���/88���n4���+{6f���u gȁ;�%'}P�H�gA,�@k/�k��M兒�,ӕ���[��$@r� �L_e� mЧ]6�Z ���7�o��0��3�ћ��#�|>i�r���w�h����ܓ֚��( F���`0^�xrPB} O���_�F��{TT��r8�9Ź�õjd�rC�!������zt��I9����0����q�*��l����	�����֫X���^ȥ��v�	]F@�)<n���o��e��Ƕ'��$@c���]!���왂/D~�4_K2��ND�g�(xT=���$�X_�u�yg���473�d
��z��y����1U\���o���w��/���J:\����j�Å���g�=~�s�2+9�{0��j�q�ѐH��=��GH[z���NoK��Y#qZH�
W�-x��l�pM5_[����.���y�5�e�ʚ��8g��*�o>����H�_z}T������t��¡$��4���0Cc"���Jϛ��x�ž�==5>A���ٿ�N���_k{�'מ;�l�m��JO ��f�g�ĄI5q�sl��1l����*��b<�
��	���)<.�7�5`��4��	/��MUJr_lb�(�&_���M�n���:��Jw)��M��&H)��S�+�?���7�@�Ǻ��tK�B��/��s����CG {����[��ӻ�*<�*��	o"x�VŰ��P9"��ϳs,�6��ϖ������ւ�k���S�H�C��C��]L�]� *��f�t�H�?�BO���{�ēǵ�t��^c��/<FG�������}�\׋�'4��s@w������<��<*����l��r