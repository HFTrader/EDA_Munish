XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-՜R��?�sk���80r#�6��d�{��3��^$;�H �$�w�t�}!��#�\��Π&�[���CBo��l�K�hʼǈ�nn��g7d����_�bvX�������o���iԫr-PkTEwo�<��J��T��NQ�Y�*K�����=��0�l��"�(5���:�&����@����S�w�9��ܟlsu���6�F_���ύU�	!'U�����ep9?G���QLqc%�̡+#+��S1ܯNS`�)s#)Vm�U�Rp��@E�bQcƜ._�h�K�yBY���XH�0%�1��MlJ�/�*�;nAw%�^�I����Pl�y���؈���ǖ$2'j+�����pGM�O�Uzn�]����{+~&�u�~�9F�Hr��t�����Z��B5"���6w���wH���l���`��:F$�zZ[�N�gtqӉ�B�f|�\4�&���1;�G*�����ً��Z"G�K5�����$eq������h�x��N��o��9*��zW �"l�y3^w�����Y��Ex�����-������᫸>�d�Ǧ�����-/Kp�Cα�'7�w�
� ��	�0Şͺ�O������6����ާb|��EKd�w����gb���5�R��6
".ߑ��h� 5Z ܩ͊� \�;��$��Gm��S`2�
`,���71tr�2,x� �����R�/i�0QP�ā�3_h���5�3��TR}#�3�n������n�XlxVHYEB    fa00    28d0��O�MD����z���0kyf��{��k�S�Zk�w���ITaG�ixBF6��so��_˷����/;n��LJ�
յ��o�l�?5;�kU�^��|���l�r�oZx�.IO����%��+�������M{ Z䂁CѼ@�U6�~�L��e!�Rtlʉ���W#j��Ozv8@��z�ʬ�^)��#��x������³�n4�u���K�#9>� aW��җ�Ǵ?�vPr����黝8�{خ����P��)�
ϗ�P�����T6��h{��Y��T�#9=5��2���Ti��~��*�T�l�hʍ�q��[l;P���F�x��9���
wc/�@�|-Y��_��9��xi�Gc|����C�͍e�	N� ښ��[7�$.��m%-D?CjO�m�hr.�C"���돲+�y-V�*֑s�L���nzD���J���$�4���`�IyV|dml7ߓ�]I�&h�!�4�\��!⏙�ͼ�b̂2[�lt�Ã<f��z&��v�ΧbgR�k��9�"-�7c�.p���:��y�d2<���M�?��O����N[5MW��a
/���J�g���O��'��atH���Y�$��D��Z��w����b�C���aq���������\�i�v*F�uQl�ᇲ�#6���c)$�#��#+;�k��L<Ot7ޮ�?�EQ�Ǫ�@ʱ,� �cf0�V�����8隩�PL5xa���u��`t�)�g��f>jA3;Z�En� �!@��P���V�X��� c�^/��`�LaoAJ���q{m��Ya���7Y���TU�ڛp�;1�b���|
� Q�&KX(��zG�Bo������Q���d96�?�����G`2�'�rۖ��F��Ri��ޠ����y*�����ץ�%��ڣ\��qO.���$8����I�nvZ��؏��i, }{\b�e���pΩ^-���C-���8�)+ �˜ٴ�>cPƒj��>	�S��K8��0.T�X��A�{��hD6���t9=�WM�q�qВK� ����.��Cj�Æ��H�Wk����ƙ���Ԅ��^w�u�
��γ���fI(���nRn,��'bb����0�f�'�M)��Ƙ
�L��M�q��XSk7�|������/����K������U��K��|Q����ﭘo��L�])��Ȼ��gaf�]�����y�c�8��Ͽ�c����4��͂��[�o��ۂd�T���-����5TԱ$�����ӵ�y2���)04L)0%��W���{�~��B�qL�]{���$��z%"�jN:��:�m��G��8���{�����[GW�����>B���v�p�(�h�aG�k#&���n"a��4S���̋�埮�ٿ#:��6�c�vJ}���S'��אUL�t;`h�ЯF{ 1�'�>������f�O�6��j��8�P�qf&ǍP7z��3Y�?��)��i�fXsJ�N�k˃��VWQE��Tʶ�z��|�+��{����=93o���u�M`�]�k�%�W�I�Z3�O��(z�<Ƈ�C6�h;��������ƯO (�v�(�*L�]�vZ���1��P9�=E1 �Ռ��(��ǜn�!~g�
���x(�3��7��lN؎�;�c}@>r"���ipN�5�.vU�U���!W�~jf̞T�k��a�>��s�T������o_~2�{eE��+�%!2a����,����X���8+W�� @(�H#��s12���v���
�{[D����p=���o#Q�*�9�.)/�3EL�]F��b��t��AP�����C0S�iTI�� ��r`��)�RW�u��p�{�IQf��2ݮ麙������<��k�����\�(�e ɿ�Ň�U>a�Z�&{�i��扠�CEʓ��t_���B�0a�pETZ�>}N=�6��#]��Qe��4
���U�X=�g�=��ZЮ9ڻ�C�7�{��%�������=�6_��P�]����(��"t	0 �����NG�䪊�P�9Bl8o��8�!���-��M�Ԥ���l�ŵb���_���*V� Gy�S&��&�\|� ��o]�|�G4S�Ml��_^���vغv��a8�^�x5��3�g²s�
���A���l�fgf%�5�6r����~��LD�N�[8<�
���~\��Ð���x���0	���$H�N\SV��Pʕ3r��[�-�_7d0]�Zj�D0��Q<�Wn)T��)��Xm�TP��5���=��&��[r���x0�!��I�����T!�@����z=�V�J�@�A4��5ԡ)H�P&y���{�B��̡���aW�[��~pL������[�˘�&�kn��#k�I�H2RA��i' G"G�d jH���&���
!�ַ��A�/FI���ͷ࣊��B�F�:�'2~��W��X�cW'�M���!+I�E�!X�[R<��f��iЇVw���"��3}k�qkI7(��k�#]�d�q�����"z��!�#�  ,�-E���w��ʕ�1<����@��ߩ��j���� �r�ԍ��aH\�kP�a��O��H����6AD_��H�*u��c�`<��74��w����=;ʘ�O �0efB<wWW���>� ̼Ɣ�7�-Z��T��LS�Nb>�g�c9Z��o\�~��&��&�����
�cp4����/+c���9���A��\�~;��F .�҄Κ�E��P��E#�H8�����"��D��'q���&�S�#�����|�l���y���ͧ� �mm|%D���`�u��*g����Vm*j���f0�IZ,�`����P?���V��*�ѧ�Xޝ����<�X��}yG�����D�C��毦��j��6['�����7�s[���~]/w��ʼ�2�l��v�}�Lc۶w����Qث��Pu����蕉��?�@�Ӧ�:o�c^	&��w�����a�{��m�M8�����@��"6��̖r螅��Lj0q`Lt���=��ߚw����
Ba����_�@.)$� �����-��'�XR�i��3vi�j�ÜP�^�EN���aY��xy	RKk�qi<���fܯgK�[�����iб��L�j
T��k`���}Mcd���M�B*=����z�iXP��O\+n���̑��c��@��"�d�v�@!:���yN(�[3�U#�@��.�9Z�Wr��Q�QF�־>�Q�!0F�'���J[��TW�$���,�ncS(M2&�y�6�^�@�&�L����k��f~nwr�����8m����8͗�BH�Ӑ/7Lz�3�*@���E��<i�v�;F|=@n��8I-���
��E�U.ht�o�>N�������#����6w�ˋ�퓩�'�6��	�l{�g7�cH��`C�甆��FaAi�e���J�,�N>tpݗ-͊��A{\-O���UA�Y�u��RF}3�M>�e�����.���/�`������x�Pi���d�wCI A��a���X�K�CQ�'I��T��oM�T��4�_��������q�gݣk�	���}SWo�ݛ��fUKp;�i�I���<Ig��@�l��ДS�Q����+�W�V�jv���Z� �(�.@��`�<dz#`C�zQ۹��E�!_��\�׶@TϭuL��r�C/M.�$�
=��{.A�X܆��T��d��rõ�2����(fYpW�Z\ib���W�6�;�\�b��K�� \�r�s� �q��&�]��9��5#�=�k���>�N]��x��H�6��	R󓵟󚴅^��rz�.�ζ�����Y�&W��ڪ��/��9��#W9�7: ��q�j�N��Ӏ� ա�ĩɳE�r���T�lU� �$�>�����Y�R��@x9��k��R�7�5,��'����j�X�VeK��0P�AS����-<��v�cl��2&F�|՜��qu�H�c�%�,�B��*�@։u0�K�޾]{Q,����?�<�%9����$4�&��+hŔ��㮋u��)�x�Yn!^#<���O�%!�~	�%{���/��=�t�F,��+Z�0���i@���^5�M(�����L�5�+�-"v/ʯi�:�a ؔ-{z�c��w y�ћ[�Z�Fϵ�#�oE���YE�m��څ�Z��i�#�N���C�F��XJ	���I8A W�RQ݈$�ts	���-%����bd��$�,���^I��Ť��H�1��yĬ��k��`Ѩ�E�b�hs?�T��~1sqȱ!TZ�3��p�<���p���9��6{�'_�Y��0�?{����0�C��@��j!��J��tg)��e�G�@�� ]Rc���W�i������ޣ{�7�[�����\Z�0��ڷ�w0�S�E�^�l�ߞ�V�{ohTQ{�����t���U���l���yi�d��҂���7�w�8��<.!7c'鞉3���bwG��I�x9�NҺg����p�4%�U ���b���2x��۳�ǿ�2y�������c�0sxF^3��{Y*V�5x��#�o�ΎSZ�o�4�O�]��yIL��n)���E�[�Iu
���<Njܿl����V�M�����ъ��oO/��L�Q� �P2�\�wb]!Y��Jq���*[Xߤ����{W��3�o���u����v�Q�?%yNq�Ɩ0ʵ�u�Fʃ�3�k.b�\�o��B8H���E~MMk5{d6&�+�:1Ѝ��Zz�욨7�P\��P�], ��NE-�;nj%�<Mg�1V���T7��oƅ7({/2я\`�Jm���"LV�k0���vd�M����3�|��@b�R4��=^�sT�M��@~�}��9��%C$Q�JΧQ�<�Y>qQIN����]f�g��?�����Xu���j՗�f�cK�DI��%��fEM���#	����]<�"�ˊ����q�8.�Tp�Mː��	J R���T�F�s�Bqd�~�p%(-L?�xRf"��.�?�v\3�{h��P��+T��q�����dNM�y%=���c��O���sm.4׌�d4�5���*�N΂���o�Q���o��4�#�S"�P�1�u�9�����å#�������(�:&fz�t�r|��ec�82%���xIV��gh\�T������_*��5�Q�j5/R�A�jN�lu?w! ��?S䡳/L�%��o��*��Bu����q<�[����`m��ʑk?F��@%e<Sނ��6=PEc1�M�b��IԔM_�b����w
�(��Sh����i��.˛	��4��Zh:Y� ��X��x����)I��Z�����I6�G�2 ��S��n~�tN6n�Ij�S�`:nNY���.L�#��W�|�����C�˽5Fu&Y�N���-G<X<�\�5�P�$�� 8�M�Ⱦ|���M'�# qSu%{-EO����ya��U��9I�ʬYPͅ�(a���v�> =:����y��2� �`�6
�-�䙂��n�ȸ�7����-mtWu���X�iT5w���Z�� �Ò���"d�����Z���Sq*�}�<�6��*O=asDu��I[���殥��%1�!�P��g����[q�8~6�I�}�(��L�;�JW�Y�.�{|�w~�WUZ��Y���uJ�y��ρ;���X�>߸b_�r<t��T4���r��
���3�1���#�9��+gȬh?�  �Y@=���Y�:��O1u�-��.�s���(�	��|�)�-)BI���Ty���q�d5�Ơ3�ƿfNN��l�aU���.आ�E��O��&�QY��i:9�p0�i��AD�!m�%����A	1<�#���)'[�΀q�� ���>�@��5���G��3v����-��I�����@gE�5͝=�=
�<<Wc�V���K8��)��u�;�S�p��9(P�R`��i_P�y��K���)S
z�tw�0�1.�$3�<Z�:���E�-�ls]����OZ�S!���:X���wF��v���>�L��).�ٰ��:ܜ�/�Zy��F��f��Xm�p$@ޜCʕo[��p��A��٩�&��q�Lȃ�l�"�����zC
y�O�1�l��%(v�7�cM�h�'6n�'��G�`,�E���2��}<���}`�\��.)���+�hT��HfJ�w��XVX�/��3'���w�8�i��q}6�׀ ��bk�'(�M=�
�*����׶P�Gw�v���#�9r���m�r�M�����T�z�Z��Cj]v��O_��7���NE@_��� m��KH�8�=����M���2�o@˝T�]�CK������|��&��h���^������� �&�<�h;�b���03)C�	������������]��	e2�}��CIE���:2S��"�'�>ˌ�����p���<��As)?>W��r�Q��^�w<B�ٽG+;\���0F��ߨ�4�,��,`k͸��Z���r�~O�t:<f��/L��R4^UI��Q�[�O!ր%�-{=1��LVm���*̬Nk*4*��x�r��Ė�dzޥP-JQء/�*ȟ^��,0mh�ǽ"�����Ú��l��C��쮭����Q��w�O����=`	h'[��:�i&
q۩)s����3��y�/{y�:��b�t:�8����>�H������	T��Y�|�����˘���V����/�{���ww։��jl�T}f� �Ȯ	U`�Y���gv���Yت\�� ������/2kp�@���P�Gӂ��,63N��g,��(��w��s<<<�"��Ih}��#{}ۜÓ��J׹�\�q5`�V����>�� �4�6�.�*� =������E������?�,jJm��+;1�P�qI}��5�]ó̊�t��Pܧzn[��i�'0ʯ�5���M��_��������"��q�s��w���_�=>��F�P	+b�Y-٪�.�R~����	��K ��)��wm@�n`{��D}��4��_�l�Y/qD3��Sp\����i�x��ȫ�8r7d+���ۏ'����y#8 �g�����-$KLՋ8>��(��}�1�O�l��.��Z@{[D��/o��sg6,�� GM�8Rq<޳�`�V�*Fz<9�-���p//V��W�n�]��)�I�հ۵�v}��� ����qD�\����e*�i�ĝ�,'�g)��a�F�h�abeF�_�S����D����"Meah<)@�VK��.���3��gT�����5]szgJa����p�w�l����`
벼�+�!���-cgġ	�/<]1}�AI dTh1��a�t{�}����훸�=}�ZҰ;����L�&`�`�Lw�d7"x����.5���R�_L�Ɛp�"�U�7� �`��?r�~9�J����O��c���ɘ�|���3E�L!����b�l��ǜ��{č�*���pi$ �k��L��M}<�=@�R�<���|�ٸ��Y�.�-�s^��E;H�ӄ{�uW�Ύ��H�o6	�Y�q�fn'�ryC��n�Ҿfg}���uf��+8թ�/Q�p�F��a,��̙^FF#2�l���� �����ЫTk�\�ܷ��%�n��<v��*�8��94�+B�-*�����˓*���A�[�C~�u��x�d�tя��_{R	j�y���)�����_� �c'�F�൘�6<2\��_�">�!���'����'�|��<��6�� �R9��x��N�N*�~��TVۀ�X�6��qT��`�c	�q�k
ƫ!�e3��)���@s��uK$j_2C�&���tU���y��ޫ��K�ڪZ�[�桞���e<���S4���<��I���򳬅0G6E�1^��O
*���9��ۂ�IX��.�l"���{A�����:D�pN�\�O^	Ж>F��t���g��X	�B!�%f�[ʂ�٢�諱6e����-�؅�Al��LH5W.behz)7PU�D��$alA���r�|G����lׇ&�a�&�t��v�R��YE�;uR�n>�m}�8�@����ňt7-��C�`{��l�B(U,O��0.�=�J�Dk6�ʻo���S_��օR��v��/�F��NOa���pE�����0�*�����B���a��&��+]P� i�ŤٲB���k'ְ��sd��?B�WU�n�W�o�>����E�E�Z"�ET�Fsa$��݇�m� �|&�䟵�T1��1�/yf��}����3�Qmo}�Pi��l��H����[3��<�
��x�5cǙ=�`h�j�hr�:�=ǣt����N����RS�FO<�q����nA�>� �D�@Lf�y��B�o+f�H��!�����EL��9 �CF�,������Q}C��Xu;�Վ�y/>8��
9hlh�f�y��%Zx��o&ς�����;�8}O�5K���k�~Wؔ�8l`Ii]��H�	���Ͳӡ�����$���r�����@&��ug�zs���{��s��7lP��-N���(��T7�%fU��m�4�?�7 :�;�$�Y��l����_�)�f`���~ZA
�[5O�~%�*L�Y�s1��Sd�-CQ�� �Ӥ�ܚ�|�� ������󷦚p�(�Ps�Q���@�E�$��������7��1����� �g
#`�\�O�C�Uq	j{)���
��#��!�h�0���MxW}ڹ>�����
�$�Wҭ�/t�U�v����o8g�uF��<��<�'U-ۧV!�Mz�u��u�q�8
��"�!̵�
~4�T��Tb��d:�9?R_�݄������ȡ�G�Fr����g�C|�`�ʚ�:���}��r�D�	��UЖ3��a��^�6��� g_O#��%��	�6/�b�.$��8�{"�+#�J�2ܲ��l원�q83�� P�$�w��+,�μ��o�.Ҵ�6A�G�B��uʹ9���w�~���L'r�//Bو���P ��K���,��iPU�4��Ez����\$�{�Y	��V�(�ۿ��v���+b�H<��j��x��6������g�e�W��s��ڞSG[^[�B�T��]� i(D�EiJ87�6V"/��w�C��	�݅ÌCG*���B<�~�{�7$�(�c���.������[j �w����Qf�hI]�2���9�+eƓ��r�Nf�>��0c�d��t4��$Hp�%j$�5M�M�p/GB>�Yf.>3�t���~�׿iJF�J��Jy\��-���9p�@��z��	j��������=�{ޘ��9�>�U�c���uڨ��g_G��[�8�����u}��y�����6< �%&˰GR��e"�������`I��W �#��p
Y*8��6f�)N�K=�x4���P���y�3-������F�A��!���b9� Љɥ�^��S�2VN���O�
_����	G=E(�d�G+��8�} {��b�h�{rwj꬝s���J=��w5��G0��~K�#�k�?�R��;��[�,���[�@a��f/N�s��		�[:�@4����ۡ0_�J��\!S�����3.m�-OğC���2�y��+݉��Z��8<�9iK�
��3^�R�3��]Q�`����O_�5�o���;�0�H45W�>��o�x/�!N���YS.�-!�{t0��V�'Q7O�	���↳�#Z�F��S&�3�}��+�V߆&���FƐ"M��l�+��A7$�8*�ݭF�ФC�EXuĐ��t#���,�{�<�[gE��Sr���x����b��eU�ˍ'X�A��k.S�6�=�`�ћ�aY��l�I���J�q������t�����d�H�Ah$�����C�%���o��T�m�TZ�y0��)����(%�	���Y>��J�V�U��s�ʉ�~ *� ��>,�����=5ج�;���F �#��j�9����x�fƞM�G<{#�-��-7Ƃ�Ѣf�J�j�"Yd�|(&���Wx;e~��"`�n�>��?�C(�W�C��<�M.��~K"�k�<ʴ����{9t���%p�{k�yGO�������� ��;��c&1۳\��7f8y������<PJ�p��n���8Ȥ@����]d0��D�8�pې
^��NXlxVHYEB    76e3    15a0�/A��0@�V��n�1�O��2_��2s$�)��o�V�̭��׭<|�j?�!8���b��z���Zȳ��W7�
��p���Y��钊��yA�[��y|��@o�΂l;�?/�`RXmh���6ڤ��*'�k��  in�b)J��k0��l��H��JvD�-/��a,5�ˎ= �<1�o^Z�>�'��ɽ�(l�����Q�R����N��b/+�+~@!|��d$�:6Xg�t^�q]���@t��:K�<XpĎ��"��l��c�xB:�&�E��<#\����"��#_��mPlA�N��s�'��5u���E�{�>�ɣY�&bL<H��r�o,-�[��;�_����N�2��^V�?d]���p�Y�InpZ�O�θf> �i��v�Ƀ����� ���~1AM��FT̿��,���0p�z����Z��|i��3M���6DZkNg�-���
U��"�{�cg�-?,)��k�x��+��)�h�pƀ�:�����z�=E�!���&X�:�*G�_�!4��a#��<:�{��K���p�Nh{d�Ǌ�_R]*����h".%	~XTg��v�fS���p��f!�_*����'�qa'ׅ��mыh���8�Ykں���O�@.����s5�L����guJ����X$�	y��kr����jT/�r��#�e�7������7��{t朙|���9A>~p�	~�g�}��3`���2�c��g�5\�6�?�s�4TW��Ȳ�a
}�`� a�s��vMX�ڌ��{v�H&��4�ZPA��/�)�Hٮ�@x���Ssh�eO1�u&���G��S�s�1=�<���u��~~`)H�Z����ܵq.Y�Ƙz�'���ܤY��a�����*�?���h��f|���*��5�C*z��[��:�F{~-wDh�\u8�����!-�w��0����ZNj� ����ڸ�e�Nv�>�!��O��F~����e"��������'�������ȀH�V�r��)]J/�+����->W_�j�S�}������ڠ ����w�A�x����A��=B�K�tk�f��2^|QoJga|�`� �Ҷ���E��&��p|�zG��R��\\'j|��Fl��x:%�ml7��Zu��#u>�rt��sq�*{o�WZ��z��U�*v%�=��{���}���uw��kg��BNIĆ�l�-��tK�+�V7���;e�w�jPy�^&���>u�ە+��r�ǥID�8d`ξ�����l�6P��!�����()]�q��®�շ�{6�3y����&��SS�BS���#�#�I�XX*�<[������S�rn<,$"CP�A���ߨ�����c�H�l)�T���e-��0
�L�U�	����(v�X]���.x����C=o[��(a�*�䝼�y�Yٴ�X�?�d���赉��) 	p!]1�IȞ0�dk��xz� 䠍bpu�#>hB�:,�/��g.����'e-�F�)FU��0��n�+� ���P��_���3%�g��&�hgZ���o��>��әD����RO��~H��J��>�&~ي�B��Mm�#��*B��LU+t<��6�r:dV��䀤���\E��]G�{eM�볁10�+(K~7��?xy�I�L�$� 
�"��d>��જ�B�Z��lZ��$X�n�-��D8�w�h���������[Oo]��P��S���e�1ベ�'��k"�0�l�`��@8m`k�x��)�kL�N����5	��6�7�*M��H��K$����s�w�?_Dz����!�x|J���&â2�KZ���@��?.��@�E���-��sm�Lig=&G����a6��[ҭ�άy�H<Sh�ѝm��C�K��.��2K=��c�dp�Mޭi6��x��2��G�܃��r��,��xu�	�I$TA�<�m������/��m!m���8�V�c<����Cl�{��"'nJ�9+]s�C�>��+[��)��[�	�"]��qɟ�(�6��@�M3���jE��_�T����>�}�ܰ	��5��;�U�M���K
�M�4"�߳CZ)��$f��M`�ڊpu�a�6+N��׻B�E�@���YD�KN��E�Q�MY5T��0��/n]�hA�p�^���&�Ӟ�iW|m}`�2S[�{����J���M���D�C����<G<X-
���:\�!�����}�Ɯ.�i�q�I��dJ�#8������N���t�Tc���x����ߺ{�����f�=%��1D�w�)�߭Ru���+yL�F\�����c��X�9w��)?l"Zw�\��+�pl+��l(��=;�EV��=^/s��]�D{��DZ�2BZG��"�e�4�Q���l��5���B�
��|)�sFH����1�i�%�ޛ=;*�X)�yn�h����
�|�id.A��?�ؕj$�c�t�BT���x�K-BN�V���|�B��/c�� _Dr((b9��`����D6�z)�2�3���E/3]�`q�F;��ZC#ub�dZ�e���;T�F!(�s�M�M整��-�Lد�q��R�N��-���p�fM sWGU����fc(,��ʒ���;�����p�u�v��l���n$�4>�CkCD�͠#�<W��{�RW�Տ���O8B�	Ց=�[���`�YFic�~���hߍ;j�r�2�`�xփJ��aLW�icw>���/�3K0��e��-�� �,��^9w��o<5	��)�`�.[c)*st��om�	�W��n���vEFL��񯠃"��0B/֔������3�0Ī	K�+�N����>��Q7�X��Z3�����"�h��.'���4l�n)ҧG� M�����s�#�PF�t��F�d�n���������z13��]���n�T�ɍ�A����Y��`Õ,e�!�huN_܇�z�F�d���d���)acg���mV���h��B��4�΢}�A���ono��,U�ȗ^^�9@�|9@��X��C��)&`-����P��uj�i
�=?�	��W͈)Xx9�?U��7\��h�� �y�Z_yş�,R�J	��t�ki,�Q~�e�lI��'��4�U[=�g��n���t=�&e����ƾ�krݐ '�d�A�f�N
ZQ�3��jV!�u"3BU�r�Ή��+�xLm��i\��1.q&K ��}/:N�	��R�D�qK	����[��>�U�L2�N�3���Y �󈦥b��G�7�y�g-E
(*qO��U�v�i��9�{/2[����T`=�[iV���i��,о�
}�k�%��g�J��I!�ډ�]&�)ױ�c�1N�J��Dzi��*<i\X@)}{e1�?[U��aOn}��T�se��Gz_�z�ĩ�6���1�|�JKjY�hza�G��v��@�{r_T��&-�	ߣ��o��9�Ҕ���6ɵX+_T+����ē)���"�)ǭ�»p��0��5�Ѵ�|&8U�����^q�4������	�Z��J���vV�[������%�n���7񏺷sJ��i^����[�Eq(H[Y���H`o�ZґS1Ӧ�C4�Mh���f��$	L-|E�QT�ػ1��w~I�Bڑ}�����nZgr�D{�>8�,'�2����O.�ݑ��"cbI���*�֪qQXO�w��u6*�����t���f˝6����D�7M��:|�u���eΞ�CZ-����3�Q+���P�[嘴&��?�$���5�q8hk�5n�L�AL,D���g��#Ef�
����`���+�WD�!,9DY����}�1ZS1x��`��g�J^N���o���ĳ���1��'�h��%(��г�MR��}P���@�DX��wq:��1��2[~'ͩM�d�<���#k�hK{=�U�{

��e��\�1�.d�H�ttæ{|��vC��;RA#�l�}�����Z�L3]Z
ћK����Sp�Y��wi��q���@��z�j�Gq�I#y@#H���$&wV_[B�ˆ(��&i�10�%���,E-|�6#�<a2<_����$>��b�vɯ�_�k0�6/Ѷ��K ,5��wJ>(�$U�e��s���F��B>K0jd!V����a?&l�Bmr\N[
N��.�������c5�ݠ��ﮇњ��}�{T��#�bD:~�ܡ/]:_f+;�V�rH���	^Q��'�US^0��Ji	В��

zA~6��G����/f�(�lv���v���o�Z���&?�V+��߽�T��#��i����rx3�UU�Ǧ=�]��ͪ�#u�p��=����7!� �k��&#�l%Km*O��+�Ҵ����Y6�utkd)����]����(��  ۓ�uwc�߬`"��X���,w� �����;`2ꐞ���t���[5�hȩ������Xc����]���\9O�yPl��ȳip�*1c5꧊�|��p	!�C�
S@���xvXB���b_��ѲM>e`YC$;M5b�ؙ7��rB�
�;J���E�{*l�6���X�'�l���l�}Y�����1�o&�d��ђ�˪i��Ǻ��9��KS�ڋ�)�]JAd�
 ���6ӸAj�F��Хa���&�d�P�S�7Dё&{~%�Ai�0e��[h�-��+!�()ڤ�k�|%9�Ē��{�ivS�p��V��l��~�k���s��{l�֑6c]��#��6��C�����n}*�/���E�D�-��P�bqBVAH��|8��i���X�V�A�����\En�ij��`��f��lPJ��/����W�J�Kp�MW/�;�RU�D{�x֊�U�?���{���a^����*4�_�3y�!m<��;l�{�ێmz0��\����(��ɱ\���՗����F�ALt��H��X��9�)��Dε*~�Tn]�݃g7F�T����.d�0��>�o��ڰ�#�/l��Kà�0~�����Up-����*��%ǈ����D� y*�>)UE��~�S����L���ȧʴ&k��+v~��=��a��[�8ܓ�25�/�̔�-o�|���gj�qIҚ���'>��!b���9�j��2�T^�.x�
�������P̓g�jź+�)�l�'FK	C4{c�>͛�@�n;zQV<���v^O�o�#T�3=y�u,>�T�mmUR�F�ǼL�[�[����0�����f�+���;���1�i5m^D)�׸��?ӊ��Mg�5p;�]�u%p �n9���J�^^�Nv�FO�/|�<)���,n�9�"�\��a�/nmb@'nK��p_��s]lW�^�Z�5+�p1�(U��A���g/� uƶ:J12��uӢOS=־;z������|�i��R���1���ڡH���0�S�R����^!s��^�5�:Ir��%X�kXuO�7�uq>�}s:
I��q