XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ƕ�&�a�$��{7�3�t,��&2>�t0�3]������ךЄ�%��[������r�p�%k�NbLe���Hᭂ��.���½xR-T�#9o!�z�-
k�I�@��l��kX��"f��ޜ]�$4�C�c��RjֵO����&Yojb�rIsf�Όil,�y�b+-����4H��C�y��L �ɫ�J=���5�}r������h�.3*9��]'�j���>܅w��e�޾[���t�>�$�C=,� �1LN�к��#��������4���e���X�p	f,��=�4!SJ:0 ��)����w�����c�D�(���T����>���HÖ�����BU����9�Kd��I���}*�.q44�ڌS����!-�x��_NFҶ��Ġ�٫�<���׾nw�C�2z|�8⭥�6Rg�48" N����=V#x$�sh
X!�zN�̬˯tCi�<v�{E��8)�*��Jr�!��0�<�1��A&��X5�ly ���XzoC�Iռ�x��?���$��\��Y_�GG�����z<q�i�M=R��_Ũ�t���c-:s���M��@��{��Ҽ,5�vz��XP�U]㺇
���ǨH����>�J/<��I� B�w���
C�r %ٟ�W�3�S-X���i�'e>���I��n��v��)W蛌v7�i�RꈻEP��"�k8�b�o'`���KJ��.�:v;w�޲N'�����>���'�����)�N�ưcl���v�AG�XlxVHYEB    95d3    18d0�݂I-����v�ԼW�$��d*]P�ʌk�)9�����E{,j	Ľ�5��d��Ư᷍Qq����x�5> �x���u+0.r�!w��/6�f�e�|�nX�҅!J�0�x�����3h����77�Aqx��j���:;�:t��6FP^�{dȱ���e��#_t9��)2g妁(������T�/�a{�
_`���ƍv:�M�z�a�W��A9��J�\M��[|�w��d�K~'�X��1>��\>K��Z���������u��A�+�F�;�p��!����-H摴!����>VN;�	�mTBTY��sŌ�i���Ԗ��W�{~wM S`��}q?V���;��ߧ;e ���X!Ë�pR�P��@	�B��&:���-8Ѹ�p���Z�<�Ո�yҠ�f������$sO��?��ގ��	L �>܉���;��t~�(i� �_���Y�,a�ܨ�|(#|�zk�ѧ9@B����E�)xJɨӊ ��]�u_��2UD���҆�@�ʅ-�,*�o�ўs"l�	z�Cp���|�jD�C�Ӳ���r/g׷�.��.F����C�2�zU��Os�8�.B�-�����g�9,6tk=�vՀ��t7z)uz:�~+$3Rt
��\M�m�W��{L.��sA����*�����'��	vk"�`ŔTi3�P�e�~R&�����-�+�r4Q��L)�Ҽ��������4B&�` 9��⮅B?J:��)�ރ�agU� �:Q0�񍡂\o\��h�(��;�"��
6u�d�����%ѭtSa?x^9 &�Pft}6��3
�;�mQ�'j$ַj�ǉ���.�D�O;""oz�Ѵ�O��#��gσ$�&-�!t�;��q��2�T�)�|�1��#Ogw�ЙeUNW�g�Y�JJ%Q�DtG�K�r��d����8�6��SAJ�1l4c?�rND���G9}�SV�m��L�
��^���JG��~2\Oz��Op0=M�X#p,�J�a2$EG��{���Ӳ��W�l211�	ґ6hb�V��ˈ�`oL&�U��/%�c`���n�$gi�}���MÅ��*  {�+&��X�����k;��R�O�E$���5�|�o�l8*f+��`}�0�]~�x-����O0�}�=Xi`�g����)�s������G��H�l�JS�bd�)�	�(�x�[�� ��o�u�fM����sZʒ3?�`�;��on�dH�̿b�U}�nu����aqIr�ݔ��G.c8HX��f�iR`�oj2O��׍���-������FG�,�10���e��<=������o�J�����PJb�w9��[.��ɘtD�~˩Rކ����|x�^{;�$����R��ܶ(A�&0>���<EAܕ ���� D�t�1"��s����)�x*�	�����śa\g4����EJ/���&��F���b��h-_�Et8���5��v�'�W��-
mzr�}�Ey�{˟�1�v7�����P���-IQ��u�ڌW�9Q����E�o���\͜ӷ~�%�4y��(���#(�A˭��>=��Y�|��
iGq�_uֱ��<�義��5c͋�}���'�X�M�����a�Ǖxپ��R���eo��c�KE���YAq*���z�@FA:��]��*�k|���#S�#��aDM��r�:}Z�����˦~�-��D5B��3�_��&��Y��t�ʪ �fx� ��H������J�VK�R��p�egq��� �@g�L��ˤ�"��%�� �B�m*-�g.Ŕ'������� �ܡ���N���M��� `'GV|'�t �V;�ƃ��˕�Zl{:�5�<�k����f0V�E\�K���,(Ӹ�'JL�> �ن�I	�U�Cw�Ʉ֬�� ���G�[��敢a�A��=�tyl�Nf��+�~�J�}��� �|�pC�Q��9I�%R�:���1�aw�L��f��#�e��|n�]7�"�)�?+}k�4&�l����yD��D�&vy6�<sWnؿ@^�h��:/��VB���HL��B�"y�F�K��1/f�U47ـ��dp�������Jb8�����G(Gj��S���b�qC����@XԜa�ީ"|��Ϡ�d��E��@/��R��!S?vaW��^���t:ڸ����t��U��[*�+�Ds��n��rݎT���F֕iq�������
��^o���C�f��*[O��<��t��]g8��v����q�h�>��ߐ�poɭq8UB��ۊ��S_�/S���F?᛽l�mR`���|Z�̶*�\A��D����q��Y�kϥ&~u;�a�G����Tͯ��h�����Z�g,�*n�>^x�tQ
l%�)��͠���nD{-A�Ek��r�̤�]5�o|"H�a�M����>z��=���CC�� �Tu�xkslڵ��0N�;�l������hY�t��o� ���Ϳ�X4����T vf>!"������!Y�p����x��{]Z�����	{!D锞���q藡B,�I�F�i3������>���V������K�K�cb��Q�e�_>�T7�3��#B,�D����&��z��%�_������>$ǳu�6<����v����P�̺�$��E�*�`��eI�Օ�n�[�+�0&�Y|�ⴋ�'j�P��I�s�n"����k�"�}I���ƚf��F����%��]���U���Ft��B�v��|�^=�D��)m��I�;�a�u���� i�
���DטI��#FvP�G�B����0M��`���Ë�X7�Dg���VHI�r���9W�T�	�E����qd1���0n���D&q8�nG!f����r��P�����g�:�
?Pn�m��m)��m��=���|X��nf?Q��.Hģ�Xs���˽I?����Y@G�XG>�";�Z��٘�x5|)�eX�P3�`1R{B�Pi��JT�D��
V��1������er��R�!�ϐ��r�۩�2/�-*��)+/�������(
jB\�C6�c�b��~V[A�N���:+��p�Rԍ�|��*>�Sj�e�ِ�u����\��c��E����0q��:^��ʍ��d�*������I�6��`�W���R��1��o�/YD���'����^��%f�����Ԍ{�D��2��/Ii�:�S�u�B���fi����/̝�适�f�U)�3�����S#����xh��)�7� ��=MV�~k��pj�^�Sqp�lH��bZ���8*= ����KL��^�� ��X����PC��ڄ� �M����zV(��4�j�W��R�{�ȿ�y��yK��F��Z�k���G�!i�|���C	��¾`/	!g3ۺ#Ū����_�壾�E�j���?sϖ�K�N��h�
57�+|j����MggM�= g�l����c_�i��-M	
���!k)�!U��
j�����RT�Q�1�X����E��f�����9����!�Q7��X�rw��Fݣ��U�&��].t��6z��]E)��3I2V���ٝ7�� �n�� q�������TCQ�z0�:8
�+��� �x�ҾȆM������o���Mݵ��?�D��#���|�[:#A'������٬'O��c/ԉv����t��Aqܪ
�-��	t#:?�~�������M\z�	wᷴ��S쏦�{	�<�eG!��U���D��f�[+Y�M#J����t���¸�������$�j���l��)i7gς����JؾO����}�o�1XC�g��x�i))o��r�	FkOB�ua�����W������U������zp.��j�Cb��U��=��nf��N��j/���>CR�{�i�a�����d^����;a;��D�d�:���6��d�r�щ��Tj�I�I|����t@�+a�h�59(�j�˯�zT���t26hTG?��l�T(��N.`�m9,����=���+㰱� -tk3���xN<`��m#?Բ<Z�.��&2��F�/G�$���U���үZ�%����Ƣ� �@y�s�'-���װn�5&�z�T�LPqD���{g�e~�fێ2��c>4�U����HVR^���'y�c�j��?�y�n�@����d���)��.x%�>��?;�&��-t��!V�'WaNwV��΍[sO������������4`�!�����m��zhإ=�N�߬4����|jy�3�S�_�Z�J�nZ������H��Շm_��sE�}�؄�j�p��2��O�+Iy�>�
��5d��k�����=g�͝/;�Y�i��'I�ܟ�������.��vҬ׵��/��$p�@��`G뚳l��u�Bi��)Z�Ko��|�� '�ݻ��bKiX���g#5�04<�8�?���/���V�D��j>���[*P�Ƙt�M�Y{$-`���i����K��#���fi��B�RY��R�h~
�4�$hr��~��+L�.C�$�o�NI����Z�+,���;M��_,?�ݟ	��l���.}��[�<�� ���p����,E���ݐ����=R6�D�TLt[;#�{mdk{��ߟJ�ї�Yh?v�g�c�VO[�s�)��]�NR�'H�G�>w[�_	��@&���8R逫05t�ҹ�z�9�Sv����"��&��7���\�"�@�U}���	4��/b>1�I Śѡ�훅���2%���!��FocݩR�!��I +%�)|��q`��-�`���>CUA��)��.��Fx�0���x���ݑ�>�f�n��3G52�;�߇ˑ���Vn)��]�G��}��	�����/-bl	���>��CW�Wè��g;���a�� sם� �݌$t��?�6k���
�ME@��5�j�7M{G�hA$��4�`�/V�Kmd3�X4�9�2~b�&ܴ=u�,gf��ޚ��P�:�+t�ƞ�X9��Eejx�)��l*�ՙ�n�4l�uݗ��hc΋]FUo�"A��i��B̝ȏ�^Jz+�!6�=4�A̛����h��s�[o���.N��q�<I���L��m��LT�EZ~٣p���P�=��R	W��2$G�t�ܾٿ���LY,��'ݻv��óW�(�A���*1d:Y\n`�;�r$���K��-m���H�88F���i�I��6P��y��c�����z����pט43��䜱�ՀNcZZ��4Hy�U�A��%�B�㛂yF�� �Y#=9��l_<*&5oh����W�$����l���؅A�v�zq��\�f8�����k��,y_ʇ�1�G�wm-O�I-�ow1��zo'��S�7Ռs�,^n䥆+�[ u��`��EkQ��W}� Fa
�*���P��Xk��>T���OuS�+�M��7�>�DpmE!�Ua����ү�#Ni�EA�;��nO��~�T(�<�坬+�Ϧu��X*�Ul �!��*P��)���96�m:zEJ2(y�$�32o.��0_��W0������3%�)����\��΢5� "MTw?�����������;��6"l��"�7'c	(�^�w��e������:�ے3���ǡ�?E[���6��O-��S�������NQ���<d���ŃO���0��U���&eb���<;Q^�mf����%l�͖����d��h�dv��.�-��e�{��R[�#���b���X�rm�6/�wA�e�u.�%��7.�PM�ʴț�����Zl����E�F�A����k)�n��A�Q�6��GMTC�t-+(��Dh��6��A��������N���/�����<�I����ڷ�Дxݙ�@'I��>��Zz	����6�Z����#��g{k�n�1m
�
� D�Q~EL�-�*�����$�O�gM�ǝ̐�F�RG.�;���xp|�1�g���D�>S-B|�\��m9}8`�]�㕝���"�T<?� �/)�6ɶ�M2p�u���K� A�z���t���.����J�!'�T��c����B�<�WFN�C"��@�q���a�f����t \E�L�����5�B�7��`t�������x�}d#��h�w���3��Y�=wH$F�M��N�PH`����s]F��]x�c����?�V�g5?@�S��x�[?�+�����Ӫ��� ���3��Js�ڦ�'����1&��p*����qΗWM�"�q��Ĳ��p՝�ny