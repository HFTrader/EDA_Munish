XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������iO�n��7h�^�\�+���j/$̲�Yծ��s�_�.̿��-J#cV�	4�>��,��^4�����ٽ���Z�[�Q��2�,@׮)3�;�W��?ӽ�6���G�������r�킕�70�G���j޻���ĈL?�gژUh���m&#=!<�p�6����G��U��?����(*������f.�S4ڐy0f��^fL��E�ZB�ґ�صM��x�P�l���=/��:ɿ<����2�O'��ho�����R�|��~|C��@���Bf1c�9����3zl��W��H�ra�¶�@s�}"Od'3���>�V|3����2q�w�ۚ�R�K"7�K�.��|��E6l���R�yu����1j�����+:i���LO��]�������������?\+׼�}���6���0�b�J�_�sL�5���<ƙ}�m���	a�6R�x��o�;�w�ὐ�ӆX�fo�<�!�)jF����#��Xs9�G���*�ymRk(���O����*�i�	k�	7��T.�(����0��E�w��C���_F�I/��fб��h���/��ĸI�O�]�Vv0xA��S�z_"�F��/=��یy)`�:��Z�ll�{��r�����Li�
���i��XX�5$�]�3�!�1�'�fw�2'� @�M����:őgFT�KE����Jwf"�JQ$�Z!d�7|�������R<���.��P�O��t\��W�=RXlxVHYEB    5e46    1530��O��r#C��8m��f�ny�s-�����_�+t*S�(�#�� �{�]�����z���R�zz
���K(p;'#ƀكӗ��F�y�#���~}������BݫQ������¹9�5�U��N�oq��\p��'[r���u��{%��tq�za.-`@�J'޸�p��V-٢%�p,r�����W�{���Vjq�/��������R�Y�͝M��v�*h��2`�E`��L.������y������<'F��O���t=�4�3�<��,O���>���^f��4�T�w� �v�6e�n�b�t������V#�B`)�E��W�6\��A���ĕ[	(���k��/��v����s��4���(��y�r�c��F��T��Z�����f�s4l�E�@����a]3�go�A� ��(d��/��r[ů�@��JX������nhӤXeA� �9���nsIԐ�S�s�έ�N���<z�?��s>�25��X�������hza�����^�X@A����`߇Pj��������-}^�]ʏ�m澢*7�?f��=����x��d����3f쀲�~���-.���I��
M�J�FlTx�F�Yn��58ֿz�-{F��9��tM;�����L5�cY߿A����JRO�K#b���S�ض럨�k枥v&7*�":!�o"=����&%��ޢ�$@��z��W�]�Hn��琟k�dq�Y�9��I�M��^�g(IП���x����%/'ſwo��)Q�/�����E��]�D��Y�)���n�m�W&�?���n�+}T�㐘�s�/L���/���(I�y���JH�S9����4~B*g�.��������$ԯnOZ�4^·�?��&�0S�5��P�� �'hKY�K���s;�w�������֎:�f���ڗ��G��/��$}���^Ҝ��!I[�]z��z���*�i��;�m+]�[Ո��JY�>�|��E��f�$�o8~�����B6�<��:�,HW�ST��Z�a" WL�m�g�G��D�r�mŽΉ��R#�\��酸
X
5
�>�@��/��eM�a�L8�V�>$x߽l� J����+��Ihdp,7�K�r-�Nj��*��ŝ����^M��3�
��l�_�M�Z�Ӥ�_WXr�U�Ce�����a�)���i�$ۃ��*s�}����F�������;^�����P�����C_��O����D(����9l�]�sZ[BN�t��� �9ؽe�>���n��d��T�K���[�z�,�P�9�ڽ!��� �A��a�������+��p���O�j��!"���{><�a&h��>ή���l���B����kD���%O܂�,~�#�6�kW֛��<��6�E�?�\�Jv[�!̚�o��~�eE=���2�<c��d�g
"�NxDE4�lUI6/�շ'��q���ИC�Y����m6��/d̤nm\	���,�/Jix��[�q�/�u]6�]h���θ�\��?���@,�gwFP�7D>L�jB��]l���-���w����^�Q	���4�嶇�%S]�v�Y[n��u�r���\l�|sO��*G�+N��ϘvL�C����u�U�>�+��D��A�zp��>�p����z��m�+��E)˶�s? N>�*�3���&Ňm�q��z[�Y�z��o�]���e�s�>?��+�|s7�ю}6�5V�� |j�#��B�
\�0÷}x�@c�/e}��1g����|�bw�Y� �*?T�¬>e'�#u��S��o�>*}0b~��&�;&�w�Y$�R��a�3ս��k^ ^�
}�ډ0�Cԫ3�߻G�(������)�̓�KP��� ������I���ǆ�����u�?ߦʕ�a����19��[;��z:��dm�-��ݶ�
�p�v�R$��4����{yCb�c۹�%����)�uX��z���[]ʿ=��Y4�9j�݂v����9�����PBr��/��0�)BI�Ulbo�a��*�%=�4A��JY`�j@J��p����Q����72��^�
��z�M����;����6�r��<.j%l�!#DQKj*T�L�p?�h�ߡ�.�R�f��RG�2<a܁�2@ĸd�eՑ�{�£em�&ՐDC�X����Y����4}�%��b���%�T�,B�̓;c�a^T�HMW?�����m��op� �{���K�Z�����g7�W���t�8�(ֺX ���٥2�Rъ;c�� �����"�/�Cc��υ6�:D��6�m�xn��p��2�ݩ1?��L��JS�.h�\[F�Rc5�'Վ���4\��UV�z�;���P�|��"BQ��h*>4'��I�(���ٔf�b�w����0��:])�%r/y)ZYtI�+yi����3k�3�.m��3;.�	�M�ک��;	���
ߞ=�+o)�MÄ�����˯��S21ͪ��T&a(�9�#�@N͑7�3}{C��4�(kem�j�������j����Wѹƴ����,N����j��1n�BnTȖ�"4��n{�����:@��c��n#�S�v��M�b�J��hÔ�~�ȴ��	:�X|����0k�M��f�#Ywpr�}|k�wt�ä��ߖ�ɒ,S�E��ΐl���t�BM}!�&�
A��y����zk����*	x/�<Ys�wT�\h�
+W��B�nӴ٥�Z��{���!}��Q�u��WDU�A֌�H��#��35Ȝ.�<�7z`L�:���H��X�<�J����[�nU@��-�A!wA��UAX�iW��ia\��5.p�9*�<����R*p���j��t�r����a@xѩ��(�� �ǿO<���BVNRX��ç^�&�'KzM:!�V�6#i���xe 1�a�y8c��)�%�^i��Cn�����ӧ�:ND����2��\���
�����j��T�8 1�ӯT���"����=�!��ٹ��}mG�8�Fg�����=���~H���ȰQ��Jg���Q@y��Ϯ�j��肆(ؠI0��/�\4�!�I�s��gO��N*P�ȅ#(ƁXGx��A���+�H؎T^�Wا�U�M�����=��� ��C����b��G�7�����7�T�~����L��C��X�ϕi���*_43Z,�>�R��#6`)�)8���F<�_�Я)V�-���<I��=0���w݉�q�{wyu`vֹ�����l�¡�_����� hC��[֤^���,�^IaƺAP��D4����&ƍ!�Ԏ���PG�3	���Y�8��@�����*��p����m���:�9$�XhW��h?�U,]Y2D;,�ve�rڱ�u0��BѢ�������i�B3'��%�w�p��:\
�v}����'�o}S �PM�)����0�9KF,���YA��E�ǒa�o41���c�#K���,)�ZMo�Rݱ�����O��� ���.@h��䤐�X�&щ0^k]��>cz��2q���o�Eo|��B`"Kw���I�2���@��(W6����s"��.�x�Թ�^;F��GV-]��!�[Ɓ���aϸ�L0�ndxB�+Q��}�ٴE u,���M�m-�0�L1eN�[�F���nB5�C�k+����^�H� 5��ŨM�� 9"
�D8��|��ʣzp3+�Ӗ�BHX`�`L4L�Ȧ��|��%��߁��$n�L
QY�5LU�K���HW�\;�� �91���;�Ɔn$HI���Sp��Ew���$kXȬs[�3�S���[(�MM�D����<�d_jHW�����	���*��j�e���XGV������x(+��>.�S��@t��'$������u6;��s=��Կ~�j��C���7mo����O���S��7��������h�R��2��!��0��:$c��h���X%�Z���e?��T���� �Z�MJ��g��M/-�D]�0;_����7�Ƕp����Ub�ʰB�Ԡo<���)�e\ɐ�����n}\+�i�2��4�����[3�5�1{�*�i�]S�U,�����Oi��
ܒto�~����^���1]��h���XR���X�ىWWh)�2ø��W
�yg.�SK���<T���V��������N/���XBI|���#b{R���(cԊ6f�+%�AM�p%�� P��$�V�#���9�����	�U��1�NAh�cUz?a��	��ڬ#:駄�p�9���u���@'�*5
�TP�@��J��/W�o+�!g9}�h�����X�\�׺�	��1/$�Y�a�%�A���6Zh�[��X`��=���8l8��ȩ� ^���-˸Sgv�-T����I���>K����+(�p��e`r)� #3�3��"&\�ϐ�\�����o^�<�o�V%U" 77�Bh�V��c�S��V*�;��=u'�kN�x��L��RX�B�'瘍_�L�����~�/�w{�3�q[;*��fA�	��y�D� %���A9�
���ӥ�-���yz.�F�J��?��S;C��(L� A���������K&��|��jѹ�E�����j*�m�R(�ȑ�����F���j�,��=qQ%o�Y��&{D��sٵ�&>*�sw\1vؿ��d�r�wu/�V��N�4,�-ٷLǵ��2R���K�QE�ᔤ�R��*O�L]-������f��������W2�Ԥ��M�Q��1������O��`}��JQ`��U�ԫ��#��C���	�s�� D<m���c��#���qR
���o�C�-�_�����>�N��Ճh�k?/*oi=v��:�I0 �`��
Ct�E��ՠ�x�_���w�g����!��/��(�|_�t���\��܆��K<t��R�a���@�����.���Av#����W�����.��M��5���p��$�1�-�sy�0K��r�����~��58m�s���]%�ێ,T��,�Tt�k�Q�ac �2��cY� �k�� f7��{�)�ؽ�j��:d%��
yG�X��Z�)�t����2���"�^�qy�'C|�u� �b���s���Y�*�<	�~���8J%�lY8��UI��'��&��<i�w��_8�����|v1�B���#C�Q��~>��%�?{�<C%G3x�vƔ�ū��݇e�P�i7�.�{g�M��J\y�R�F�[I[�y��T�NO�ʸ}��Y����6!>�M�_�E��k�G�vHP��G�cD��0V�2��-A�Q