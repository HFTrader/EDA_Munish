XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��m��-)�2����Cқ�h�R:��>g�x�tP1�*��Q̉]=R�9ҭf�� �*)'c��K���9B��Z��6�}c7�ˍ4D8%8�h��|WZ����j�s[i9���)��Y����)1�e:ސ=D�ns�`&G4��J~W�o=��a��"�܍o�U�,t����8�j�[�I$hG������fN�6�oy]�2S&�\PS"N�.�R�b��o��n�����gQ�!(hH8��p*r�k�z�<��t��͑���}b���@㈠�t��kVE�.U#]��f+V�iH8�����hc+<s`٧��e��\���G���J�$k��=)ԣ��$1�Wo*�+sޟ6�$Ʌ����~�EG����v��#����Od-G0Z((��uw��ML�VH|"���e�����}7����5B�T���E�6���ĉý*�@��Z~��՗���a8��"|"F+.=�r���;sZ�Jk��k>)#d���F��t��pJ��+�F��q��0�+��\��b^�}�O�:d" �&�%K��	�oжMuG��?���c�1�|�d�=(ׯ����~b�?�^ul]�g	\�ܽ3�����n'�_D��h���
D㍒3��|m�����q������	������6I����v�e���_c����77��}1�m�1giv�D���l�^�l�ZF<dΘ2Z��S�S�R�M>����'�hAn\܍.��ӇLTQ��E@�0u�X�XlxVHYEB    838b    1770 JDA�`�}	�� o�ǿƋ��'�;�3A������V�rKӏ�r��<0�j�����vy��}�0�](	e�s�H�×\���
��E;WT~���;:��r��oĄ�M�w�����$��9�hz1I�T��\>��N�@R!��b)E�Ν!(c��.�6��#�s6��S7���`+P2.mJԯ�ÙP5 �����
�m̎-2~0thc]��c\�ڧ���#�����F�.�������Q5�9���X�}]�4�PB�<���"crn��W�|��o*i�Z�E����G����F�<��1{�$�G[ �Ƀ%�.Ȁ��/`\ϒI)�T�O�*|� ��*+�؏���Z�z�PB��<�5�b�@
m<��#�-ȹ�)*��=N�J?�+VY�,SX4&ܦ?�wM�����OTm�&�L���&�&���na,���_c`Ҹ��K��^	�h��m��x�p|H~Ԏ�c}F�UsJ��d�����Ag�_�X,�7� �yq�'�����#5��P&+x�I�g��Z[�GQzN og%���A��N�*��}��I���ې@eF�wҙ����"<��u#�^�T�$Z���_m�<�M���f��Y:��v��԰Z������Ě?+�`.ɢ�:�ޡ6�H�m��T�wy�������΀��b+K��}g�3��rE������+4�Fw����fcYe�lߔ��W�}��3ѱY'�3�#3:�]f=�ڜ�.�Z/`#�j��
�[$`�LrS �U8�������4=t/�_��rؖ�q=�A�v1'˴�@*Im���ß��B��}�ڦ����@�6jD�L��K4rۃ���¹ɘ�nn5�}�*�����p�h�&��$7�*����H!`�����5�]�O��2�6
�Ql#�R{�@�\�F9��Z"�U��M��_�v�5]!�z���c�f�*���v������G[x�ޞ�}����2�oO�E��������o$ju�}�-(}���j6I"�Tgl�uiO�>��G���X�$�}E'��ST$�J��*���d5=��J��"�����H!�[�:�8gQ�$�h0�!B"��b����(�y���!�\�F���3�>�P�Zr��%Jx1Z�c�r(���/6�)��y,�z�6�Lf� �0r&з!��	�S�u���:;>Y�`Y�P�R1|�웈�}S���Q*(���|���ҥGSd's�����Xi�ɓW	KG{��^PlV��M=>,>�т�%�jgs���(U]@���q���x~_�ehuW�G�9M�s�N�{ )�1F:���3b��׈���v�+���,t<"[�)��c֊װF#���y���gU�CA0,�[�I��
���X4\B
!͇E�a�����T����f���9��8f$�:����� i�Q5�´:K�[_����|�ewY/�F������¹�ٱ�6C6;�!阳�EU)����ul�夎6̏؅�;���P}�����Q8!�p^,�H��X�_X�XN��IZU�f_#���Jax���q9L����f�kg��3�������Bo�(g��ݪlX��Ku��q'��o���R9�r]���ӏ�=�a98�0p\%s�Ss��mz���ݍރ	�0�&�61w��2�z�A��Jᙽ�����j����&���X��;�.��;�\s$V��������&�Y�'�x����G��*,n�>rLI������Ƨ����� ���1��R�Y���Q6��"�d��McV��<v���C�"��"m�J��u�EiH��*��/
t�������.��q��Z��������$=�ӆ����k`k2߾7���T��ep�"$H.tк�y*�ϖ�N�h'*d$F��u�Bg{j��P&#��|v�s�A|i����2��+�0�@_ݽk�.+�ˤa{����:%�v%��xW�����:`x��O�v�p�K�% �� �ֳ�����Aː� y��6y�"��`��P�"]����v���#,(Է۸`�1���m�"��Ăf���4��>�b Z{E\��N�n�l����ܲ�A���d��;1�꧋}ک_{�����D����C���^:9���������?��X+�4�ټ�T�t�����ɾtP���myEw���Md�_�s���[lV3Dm�7��dW���,�Ǹ��ϐ���[qF�an$W�ǡ� C��/_\ŏ����ߪݰ�!e(&Ԏ�<*�`6dS�[p�I*�$�ng�(�71�>�����9T|���F�1�Ȓ��c �&Q屺�I׻��so�����cϠ��7�v����c��`%�$Qn�����(�d;"�4�C�D�{���\un��^!��y�����hG%����3yVB*�:^!��>�� Q��j���	��{G�p�l�g�M���Z��Bx/�]��9W�Ͻ�nU*R�;t����Aݣ�->~;ܨ�B7`{L%��#�]�j�c\m\���RY����y맼W�&�V�c���ܓrP�ek��(l/�px#�Y��p��g��F��F`MH����&ge$#����9�F{&��<����uL��L� ��Nӑ�^�FƋ���8Fح���3$دK�뷌ɜ�$���m����%ٿ�'6�r�3���3 �7���­xHX�vR��U���Wݺ;S��5s�K�~P�ns��B���N�D�hȷ{I��r��Yҽa��g�E���<����%�m��|!u�~updt��a��V���D��3�ԋ6�ꞧ�k�G�φ�Ym؊��f{=�t��=L��)l ꥝Ep�	��}[+qR�,�J�%�@�bw�nl�Gɋ��CVu����ܪ�/t����	�3��Z�C������`y���<ڹ�m|�J�|���z�ws<�(��M~���h�����[!:��Y�0�c��;2�~���i~["S;}c�t����
���gJ�6�Ǚh�� p�����$��>
�<&f&!;<A����#o��-�sd� zO,,�Pi����?�PȌ����*�8,��J�Ӈ�~}�{V�1��hB�7L�=�W��h����Ϯ�~l��$=��D٦;]�,�U�Cd��S&��uԠ�K�%�aɖ1�4h�6�2g�Q'c�G$��;�\��w���#���bԣh����ZF)��/ή6ʹ�N�SZ�~�j�a>�y�Ρ��= $iaaq�e5��L�f{� �sU:�`��� ���>��Ջ�����>�N7���,e��J�aM7gCUtg&���Fe��~)��JGL2UA\H_�����vj*a�V*o8����3"9v��(>�@�J�QЁ�Ԫ����!�C�����k�^�fJ�kO0ԣ)=" Bk�>�V��R�Dд���������i_^�m������),�$[��i��]�|�;�iv��)�&X
]�ˤD� HlE�I�ab�)�H䶹�`��>K4n_c������(�_)Ĝ�u� ^l<�����@u��gif�u�����S�"E��\Y|�lq{����6_�Qf�3�����Cc�)�-�"0Q����`�����ל�M��P�*���X�c��,��Z\^�������Q0���������b�K��r�wW{�7�0�r����_؞f���@�}�L�ȼ�Z��r^xb��<ܢ��VLԕ9:=]�$��~���A_���h����A'I#�ѱ�Z�71��P<YY~��)_��@����t��&��������7�H�§��S����	�� ���4z���^�[�����o�/h�����P��V+��=� J.I������XB"
F��h�o�ͫ��sPڛ4Z�S�k_�ƨ��:�4,����LHʎ���ܑQg�[K�5�t�	�."�Cg�B����X�oo��=�:��\E��-g�nV҅��PS�֕\�����v�\֛����-��+���n�\��	�t�jGF6E��h�]%�!�HC��o��VڄK�22�Q�QĹ6h>��G-��m?����1�"-fX��5�?�b��.�EYq`�p��Ǐ��D@7�x[u�g 9�#�B���5�<�g
�Z�	ҵ��3�������U�4Ґ��f�x��i�"���lQV~��b
�����	�ԃm�oJ����������z߉^�v�@�ҽ��ĝ3]����l�;.Cz�G�ڲg����l��(��z{jT��nN���is��^AU�������D��jYI�H�M8����i�85�W�!�/���-j�f�5�����=%\ΠQ ���DMP%ϑ�������j�vޟZ���� @��1��@� ��E�0�MJ�������p�I2�SadX֫��x���9�/]�`�I��c��v�{!��g�|V�%揓�,8�-�W֤�,#��T^w�W���i>O@+�\�m�i���J���;"�o2��x��Wl=��RN�{�p���@%�{��1RHLuk+�"�k�í�м^���k�I0�d�-�hǆD*Z���B.��uL���k�^D�`��+��ܡ��Z�Hi~�XÆ��j3MѴ;Zk)���N��T|��u}N:�x,z��5y��7���1������T�VI���sS@de-�r�Q*a�o�U�'�
��T�%�*=�ʛ�
E��S)X>B�J�|�n�f����b�~�����W��0G]�%7�HQZ ��j���Pך�W���4dy9������:^�V)ٺ�sI'bq��gK�ؐ���N���Bi�%� s��t�,��@En���:7��L�Z�	5_��'��	� ���#z�+�Oβ��q���a�k��]��3-MW]pPt,Z��:F�^Nw*��s�
h��[*�?\?�x��F��M��)-b[���JJ��������i!r�%�i��>"�G��˵�$�R�H�����?���t���`�qbV#w���jU/��Ep�-��V s�?�刯�:G�՘���m��=L�	r�"�9'�D���{ó o���ȃ
Nr�M�H�nfS&�#��#��?b��.W�`�[7z���N�YN�7�ts�vb���W�L�H">#�O��6��eƫM/�s�X0㌪G�B�A"c��'�}�-��8/4cŇ�çā
E�F��;�r�L_�4����֙��w�'�M$���.@]T��2eg=�=oS���.�B��S>(��i�q��8�焳��୫���
j�Z]o�+����(8�����L�M\Լn�-x&��ozJP����Y��Ӭ��EpO��.�LB�-�-���.V/���ʞE:��Xv�+��kA��� �S;^����^��X��h#�-�`D����UNDܹ�Ti��]�O��M^*�����L��En�8�ާ�*��}�M\.ր���`�}>"�����O�mSrU_�}g-��g��S�(���E^#-��##s�jQ {EX 9L`[K�s5l]=�!ƨ��	�XC��(V.LH4�i��ZF�D�/"kX����Rڢ���sS������H��@�k'���}��b���?O���EAȩI�N�oF�mӳ�as}l��0@1���s��ȉI����Mn���X�\�a��'���}0����&-�Xy^��9�
���t�y�c�Qzۡ�[U�}
-����b
>��q#�Z�����E�2&�޻����_��A�`�?g=i�u|<g�1a�����Qۻg���
�P�Ӯ
/�����%��+��p�3������;m����-���r�����~�Q�������=n/�Od�v����B��P��
%����y�����6Џ��E� �'1�@���v%-��;y��/��ڵ����>!i��!�(��j8ŷ��6Gg����)0d�mn�P��ϰ��Zܭ���*��Q���Iwzq�B�