XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����V7!l��8�p���O���&�zށ�L��$�y���a<�aL�,�ޣ����^�jcCP��� ad�'�ߍγ[&P�w�2Ɛ)�Z������@����~�/~fT�C�&�U�5 �� ��$�zl����0��:��	m��E����2*��gs��1/�N\r�t�@�GB/x�r�	�]�]d���8f��;�����-!&p��'ɖ���!aS��|Z�g��l (E������5]���"��X��`S��ʝ��-��t2K=͙K�Y�Z���\X����ڛ���~q�?O�7+��
sr^aZ:�+	�5fۼ|?v�!���$��a2w3��������!g�;��(o�f���W$Gs��^V���O�Ԁ�i���5��1]٨e���������>:*�Fx>��d� �ʠ��U��>�LF5��Q�S?P�%�P����}Q��-?� މ���+[^� 1�[E
8cѽ�Ir��a��\�]:^��?Uj[�o|p���b�D�� �)���0k^���/�k����}KeԥHF����
�QJ����D�@ʴG|��/�',(��o�|�1Ɍ|��UcVz+��'�3��!��?}Iq���,�f�\&lw��BKw�L�g������ypV�^0s`e�}���Tm���1�)�&r@]���������Q@�g+�=x�L�ڒ�4��xdX�I��0E�����u�&Ò7�BV�k���]YD O	��Q�@����(7��t<���N���XlxVHYEB    5909    15506��������J;��Qth�['�9������Ɋ�# �J�6m �c�q�DW�z/�[#�L�R ��eGP5��@W�x;�����BD�s:xd��f�3E�6}�R�<<R2��6�����9�F�:+'�q���&Bw�����x����іy����,V'��� ��%�M�7:�\���q=��@%Q}D�J�~�λƎL��C.���v�o�IN76���(�QLv�Jiln�1����=���"a��O��9B�-7��i�����^nM�\!A�IX�M\BU���ʋo�������V���h'�ND��m�p�����o��{`}�ia�&� �I_z�(CZ����m����a�����<l�V���_��$I�4[��F[�e����`��d�*�;�g�8�ʾ��<g�&��U�L�T[�:�F�Wi��E��'�8^iL���N�g��yu�6�}0[ew.��-l/})[ߎU!�B7#��SeP,����k�H�ܧR�S�NY�+�S�N�*D!z���q�l�4R�jZ�z�����O�m��,�sg`�@`�x�=�p�7�Y:�߄���]����88v�j���l6���
o�0ۛ��z��X�#� �`���d��w���fx��Gҽ9X��GG��~+n����V���q�[c#ۘ�4]>:ZP'������l��i� y��E�K�L�ߘ�(�kP�QahOU��D7e׾�^f�o,����De��L_ف'�9`�x~�H@V3w�N��m���.9���R\漵A� ��l=_�w�BDK�:mdN�B]���=�"P�hYӏ�م�fA�Ĝ[!jK��h����6+��~��%~V�v�˪Χ�}`V���f>��E^X�?�9����Ƭ��eg�O�?6�@�) (���d�������̘�])<�I#��	 ��M�L���+���D �l	�L�O��yޛ����TA�R�i��^k�i�:�㥔W��j���������G��*I`�J�)��Fy�o�y���s\�]s������W��YBN���2�FO���3J. &��S{KZs Ŋ< m�5�v��Kvű�O�Goa3�\�Qh���O�k�3�#b��ʉ 7(`�u_��Dɚ@�~��&���c�>05�u���f6ց�v����`��`��������}o�m��������Z�,zP��_P�[�i+Jx��l�]3r#J�F%�v#?*!���XS�� �E�TOA�h�4S�Z�E�r\NIܺ�X_&:4˂|�Tƾw�[b���u3jX��ݟw�fuU<w=\M�Dw�י��"G��Hq�A�Н2ݺ��(6��}l���d��]�Aٶ�@ja���}��J�۠���JH�o~�����70�{q�B��j� �
e8���;�5'@��P�{��ܠ���nIlб������Wh�����;4ٲ�xX����<�%�F.�����Y=V��C���.� �,Ղ�Hm��_���':q��U�pz������%����]͝������E��Gw1,�';��BI;���q�J���P̀䦲(Q����2�����N`��8�o��E�Z@�@E/�:Fo����#�:3���^�rÂB�E��vcb���\q}J�@���\۫�%"�f|�c��{� &,�ŉ;G�y����ݾU���m��uJK��J�(��ⲻ���?� i�o�Kê��Y����]�ۖW�jS�
�#��\�fu�e�C�תX�6�}�5u��ۊ��gv��DZG:w������Yy�������U�@��zU"��u�#-1{&~%���r{��� ��J��djQ}�����U.��W��c_֘Ozt�А�3�8�
�|�q\�S�P!ΦCCy�&�kތ�gp$~c���n�Y�&Ƈ�S��
��w�u Y�]�^�Wy����&��ǁ^�GP��|U��<�ǳ�A��!���G`Az"��[*T��9���}*I��Cɒ�mh� �m�� �-q�[b[6	Cs�1a0ݯ�}�`���"l�w\H�/�Vbs�LM�"���Xv`~M�E,��|�M��_t7�3z��Rm� L�چ{�}3��,�!�ip����g,rZ�@:�J���>,��0��Z��%[=5|�P�93��U�P�E�6i���~��<�)F5�37���=�ҵ���V�{���,x1���A
��Bg(�b8^���L7�z���x����~�[h��BЗSX��8��6�y�,��o`Ɍ��X�9EӮ�t��32>�>gOS4���^���}Rp�U5f<�rr��X�u󥻨b����� DU��3��D߻��yf�O�����e����vb�Ə+�C�ٿ���±fa��Vw$"�g&ps�ӊ�)��k��@Q�^ūg�!���U��Y��N]���fQZD���>L�4��;�^���J�Z����4�ϒ?�B�1A���.������X�
z��f�d��75e@�|T/�qd����z�pmq��D�$CZ{�3�S���qum��!�Ae�u����ە2�8�����K*0�z	�|wF݁XG�BӮI"�e,4%m.W��Bp�W1=>�?7��5�(��9_,�J��!b�}�/�Q�,1y��:��,	���j�*�˯�U���X��QݢՊT�幟o�Z!cbӻ�ڎ/�ީ\�~S@�j���X�0���(F.����K���i�7��#��tN�����fw!�WN���l���al����Q#_��V�5�%�ۙ?�������Z����}���b�3'��-�<F�8 �\�)<��-8p[}���ƥD���yrT��Ā+�p��>؝�꼛���ԛ&�5�U߯�%��U�ofg��7��{q_k�_���m3��L����
N2��͐�`W�6��Q��˰���������O�o�-Lɑ���D�pY��ldM��꡵�Va�cn`��׹}��ν�P$u���*"�T��C]���u��\*�		�pT�bs򇌛�Lg!sD*���y�)���k���_�6�-�S༓�?��}��3mp������@����gP���Q�@[�e F&�TQ$��v� .��R��f�5{žM���l���֫[y^�2�;�rh�Fy/=lQ���4�hժF�Gжk}Ri�ajM�*nહ��QB(G4n��A�b��?0.���_���e,8���M�����#�`��pٴ.~?��t#A��8FI�&�/�^��"x���)0�g�oV�jI)@=W0��̳�{U�M���f�PH�����Z)��S%��,����ga��o{sAn]�0�Mp/�N�)�
!gzM��;�ь���fO���U����-7�=R�"\-M�R��B���!�oR��'M+��w��>k'�H�*{|�*�B�$�1H���i~��ô��@�"�O:�V��+���ړ��c��Y��ff�z�{�3ٮɑ�T����	�Q�ȏ'���֫#�%:�aN��X8��N�|��{ť��r�:M�#���{�СT�˼��5�G�gؐS&�n~i{�I!���>��]��!X�|�#y�v�ٛ����*/����~� ��wLa�ت���5���6���qm�p������E2�ը�H�qS.���ʱ E4������/�&�R�u(���G{$%%�`���:����v�fL��0�!ld�#[���V����}�t:Fbw��53mW펬���7�Bp�-(��;C���D��R���~B�	P���'K��8��J8��9^2r�16�#��<� ���_���ݸ�V�H�>F�g�	;X�/��$,� L�w\�T��z6�>.y\1d�FZdF�,�.�@릪�t�����\؟�7����a�*�ɑ
��v���6�"+���'�/�|w�ٽ�'$���s��$�ڹv��i�Sy�5�",K_���UݑT�n���s�:�Q���K��o�H=��p?΢Y����1�_��I��i�Ex�.��c���7��H-f+X1�(_�T9)����R��6��㢇�B� :��W��RO�ꊩeX=��Q��1
齐N��� ~�)HGx�� r<7Q��̻.s��샙J0�Z����M�H�H���VC%^����#�ECݰF'�;���'����m���z�N��ީ�>w��հ�H,�[`��6�>�V_���!�l�Qo��xG�=�k?&<Z8/�����4�o0wӶ�Wp'a��35=�OU�^KZ~2ѓ
�Z��!�ʲ`�b89ӥ�&��X�YX����@�d��O��X���� �g�1����)����y�q�7Y��&�M�mL����
����s��⸱=�}� yv��:<���g�Y)xk�4O�RUk$]ۘN��ڪa������}_�K; �$V�Ĥ�/�̯'@1�k�#��AN�؇|�Z����DL����Pz����r����pa��V�03U�+Ӆ�t��F�"A�n��&+[�;�����u��i������#j椴���E�SG�YqX%U��I� �_5����7��ք�c�HB��<����8Փ2�	�ӳ��,P�|��BT,¾��څ��誎f�+��&��i ��iJi&[rP)��6t�|��g�P.�bs�rHz >aqS>��d4�g &�i0 �v3��J����o�{@\NG��cSo�44��u��lY�����Ta<�l�����z�	��B�(�|�����^, ����AGu�����?�U�o��Bf?q��=%o�f����2eq�WxhmV-h��=�%t2w\�O�m;���1������L��ߴ��Ĩ�y�^�~����ؐ���fOh_�z��{��XF��{���CA؉eɒH��QpN�Ǫ��+=ݷ��Qʹ�*'s��U�����"�+C� �6O2�e�,�
~nNx
��N���ʡ���V6�(��a:T0���s�[��cZU�Q��z�s0ib�,��Lo ��J�� �K�.#.�m��L�T8��6�0-���bA�H�*^���Cm��M�-.����S9�_^���ӫ�|G��Ѭ@槤�*�4�D��m�;���]s���اR�4��y�?���)�}�)�u(J]���+U;i�.��ĝ`�@�m>*�|��d&ʆ豠�;�����2�%��:�$j�v����K�FK����|zZ)j5���03��.���]��F8���]s��Y�����N����D��(�eX]��S�gr>>�dv�W��v/^RB]t�yR��CŜF^\@��()iE�Pa�