XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����w(a2��`L���a��n:/P)�������k��g�n� OgW%�k�Oqn�F,��5!h���:g�\"d��?�o���փ;�n��\�G}#u���͞���������)��Ae����c�!2�XJt$w\xB9ؘ��l�� �AV�&��������'vM&Kx�{�mܺ�QԓdWI��q��P4��Z�W���1���bS��o�۰��q�ӽ�tC�Ū��%j	�����_�-�����r
oUH8�_��S�Mڳd'�e�a���|X��Bk�:ȓll�:�#����B���"�q]J�Q2,��Q@���I�|�#JF�I��N�f�l3�0�xP�f|��J���S�I��ы�H�k�ׁ�|�8ܬ�v�ݬ(�P,��2�\,L��
?̳f�|<���$�2¯�Y��Hv��2�� N;��%>�dvEM� ��|p��ì	7	��XWuމ�&��l�����M�]�;'�ab \n�z�KW�P�T�)�p��~� ����R�,��W��$���2�!��B��c���x��g���ٲuQ��a6M���Y�3K,o�ί�	)�>�ހ$�4�q���W ��
/��+�.�� L��s28��� �1Q&�m;G��&��R|����S��c��~_W�J&���\��0�����!�}f�D�0f�t�%b��+�aXm3ח�%�>�����u���:����P��7lz���N��6Κ5P������]XlxVHYEB    8e9e    1d40�nvb�"(��pC���vڛ��l�I�x^��o��b���0���(v̷pX	�f)Q��N?V�Kϋ�E?�-z�D>�x�$��!o8�>̵���]��}��T�|�  a��v6]/��w�-�c��g�������ǂnPo��+w��氒Xd~�E
3�`�@�|�;5�5d�%�{����iQj�'1.��{��U�o��0f|D������N^��e*~)���o%�:�;�Z����,���N�8�1�
�'��qd���s�3��=��q@�,ɝ��+����y
Y��@��/���mF��5A�5�%����]0 ��L�^����D[GM���(:�%h����:��������i��w�G���=i�nPC�'5~�:Ĺ������퓓|� �vs���>���IG�f��S!��(L$��>is����j���f(�1Ή�g��\,�������$a��X��pn交dui�>5��/�V�Y�\�to���__G3�]B���z9�FC �(�BexS���M�Hc[>�&d(p�T!)��&'ͣ��%|$���F���e��!�=>ON˒��H�w�0���v���Pԥ����d��c5&�\�[�I:F��nH��Q~t��z���m���ǌ��!2'D���ʟ�ж�@��4�7K�r+���*]�Ƭ+���q\!�V�ˁ��r�����=�Gߍ
�H�������;�\F��W�U��h	�<�3cӄ�b���P�Bȡ�!f$ӓx�;��P�j��*	"�����i����H[�m/R!k�sk�	��[&���a���OČ���*ﴝ���j�&_N�SK����dG��h�^}T�0���Rؔ��\|
/�m�Aɋڜ��w����=��<�O��v2Kn�-�h�F���PIbV]�#c��c<��0r���� ����`��!���`�Y�C�7�G�2���߀V��+;\QM�u���g�L�{-�����m+��jڈu��Z��*jp�z�ķrv=׼���f��qK�o�����L%�i3�~>��I�tq�8<���cL?����[�����Z��0I���;Q#%.�04�>�M�#@�	��Y���v�:��IϢ|i�+V7p�F�B���U��uW%��J��^�U��ˆ�����L��H�������6�k�*p�.�C%M��3�z��?��G\~��+	�x���>�~�Ns�du�����%5����� \6�2l��+�(yc��'���(�����*��9nw)v�^����b��&5A�K�C)����c��x�J�C���w7qN̆����B��29��k��$҈���y��鶖��dw��ǔ�?ٮ���,���hAW8���]!;��4�a�_zC�#�%�7�zJ#�����I����Ad�Er�}9	�1v\�~���/�6�s,&��,(��XrZ<Wo���5Oi:Z56%��W2��3�t�,[�I*5�nF�䢅�`�v�<>�� �my*�y�����Q=E�6���T�dl��j��>���}0����:˦�y5#��q!-�'6�1�$�҈�/^/�Фy��{��a�X#�/ȸz�N�g��4���x���xoNZ�:��T�V�Bf:4��A��}Xx�j�ZJm��|Vԩ�+���6l�%M~׈� ����$����|'al�#����sޭF\hBr`��4W�T}��7�MM��M�k��mV}l*I��@ѹe��1�p;kϾ������J!�*~��cU*G��Nu��8M7@�$F׶�|��ri���������P�����0��!'�J���&�����O	��wF�/W2@��tq`���.�|tv����F�:5](j���皦՗��~�X�����%A�Q��"dvD������9/�	��8Q��L�]�"�������{3"R�,ܼF�j��Uۤo�� ���F���a�%z���Qُ�M�nҠ����|D��`so��b~��M��Z��|�Z�HCqS���&i��yg�X��1�0�r�-6����"�.^r�#�� �_JF��N��lř�Օ�x��%(��b٩�Q��	LT5�s3��=�A]��R��>�7)4M��n���&���=8���?\L�Ydhm�����gJ�`�K��`q�D���*չ	m�k����+A_�:���qI�*r6���;�/n���jL��_��E�^��Ծ���`eSk`�:��������� f�:V'��P��iJ���g��jU�%�����\<.#	�է��z�Q &Rx*>��ڂF<So�!�v =�j����^j��=5 �h��:TɌ�@~��+K�c4�*k3�����뺨�ԅ������d҉*HԳ�~��P�[��Ĉ����fKui�®0`�e�ՐtV�Sab��LAJz��ߖzKR	��t�H��H��'py"?�ԶQe.8�Z;�j��Wb@�A͡I���`�$c��Y:��d��G�"���M*;���)vi���Ǎ�>��]u_  �SE[ط����<��}gkYMxA"�d��{q��h�W�I��\8�Р�O��ɶ?iQ��YCV6۔�r�C�
���4��X=E����b^�b�/W�b%�sb�q=�n\��pԜ`el��ҵ�v"r���@�C[�6&4�$��b!n���vi�PGt~�޲����0;��_}!<Ѽ��Q ɢ%;�?�N�1�ǟ��=m\�5u]u��5��t2�y����+/	<sZ��I�J���ͦW`�5�6���o,V�=O��v-�����HMC�� �0\��!v	g>6�nu��MD�XG ���o�K��W^;��r4'�/�i������1Ĭ���>*0i��p���{� ��`Z9�تF-ٜ�5��)��|�g�Lg�Q �D�iDO�?[O+�i�|���]c\� i	����9S+}s�KiE£�i�p��WJTt�����4��	`vr�u9D��f�@;G�LW5ny���6��bO��̦i���{�&�<~ɜk�ļ:L�"��k� �� >+���ɰ�!���Jp�C�K�G�s��_��xM�"4J�����k1F�s���,���Ht��/�1w������r��@G��׆|����8ӆ�����I^��� ��m@F%vG�;-�s��.��(�O���W�t �R��
���{��8�i���5�+�|��`���d(�ȏDM�Ԧ��40����T��uq�������7n��q�L,����ʟI�b�l��?��U����m����hw�A{��d6UT�AԻs�)�����B\��q�O���;O�5��/��lCq�W�>�иx��uD�����l�TΞ�5�-2x�,�+6�ߥ����h6S?��7[���'tM��v]���7���g�>w䂔i΂��2.����V"�<��/.�W%��;!�2�(Yj���M@�q��ō��ѝ�2-������v6�JPSv_@�X�)o|m�����39ch�.mI4*6�z����tF���9ʞ�����l!S ��K,p�a��OQ�� ��F���O�V	�p�V�*�6���%�@�5��p_kǂ�k��?8VՄ C_\�m���I������vR^� �Ly�A�Xp=��W�����,�A`o���j�6�I-�'_��i0�����Un��LxBf͘	~��,��9�>I2"���Ώ5�&{6/�ڞ��J�~�Ǯi�(NBdM�Ӆ�2ulc�m �&���9��wDc&2:��s�r��.���"1>�3��۹����R=	Iû:.Ϣ�w��ޢ��&�IN;ǫ6��Y!�� {[�W�-��e��S��i�	�eй�7�0{Zf=�=\��ߡ&�/�6�β��?2�?�����v���MZ�(� ]n��T��PO�8�Kh�fͳ*���Ēe�!� ��$�3reԤq���Qڢ���vPL���fX�_��G;)���;b, �d��n�9�e�/���id�C�mcj�'O$���5˲�
XF��ޥ	����X���Y4֑���r���|-L֘�g��f��ƨ	��4���<Ȥ�ۜ� f7?��1�_I�;��S�P`���G{
>�jqu>b'�<��3>�d������_]��Ѵ���/� �"s���Y��@ 	�S}��M�c��]�ܾ����R
$6�^x��>Y�4�2r���C�ʀ�l�����m2��ȄE��+��{�N\\��VЎE�������4Ya��
w�\Щ�mx��ÆI�T��/r$@��1�bq�/oH`��<sCke���tp5�K�A�FI)�
CegXq�ƬF�°�=�8C֦�)��	 yIg|M�	��$�4ʍ����E�OlA�"�m|&ׇ4�˘b8���X�4A#��=xL::i�1�,彦�Ju�A�t��&�*l�j,��}�#-�Ud����L�mLՆ �5��sm�,`Xv"|T�D��r����To
ȡ"�+��R41l�N-�jh&��)��n�]���jGˍ\��}�q�l�2��t�/��-�c�"�ڃ[����tp��K�������ڃ��|��E���a�Wj�MG�q�Z�wȃ����!e�����&���<s��%1����fL 3�d�A0^Y侗v���[�g��d�/4B��qM`���(��1ڦ�5���O��I*����is��==\��0w��}��廆kSM�������6���O�����B�,���#ێ�X�w犏a^�&��S�A �<�$�8@� 0Ҩ�J��]�qK�<oBU��u��)N������n���m9��QG2�{��>���Ƴ6#6I?R�ƿb}/ڃ�٪q���isR �r�oKp������|3�q�%���u�L�l�l�i{W^�|ݮ�!�aR^����DW�v�@�Gͫ��Z��n�����R�P<��f��q-�	<����^�(�xH]B��lj�qP�T3Xi_hbseYa���[C�1��L{3�ϸ�y���9���T��8F���	Q�0��;>�|G|>�����$�2�?*����#�H����'��^ͼ�k80;{����w��`9�}��f�u��Z3��ؘ߁5d�5X�6��k��E6N�6�lYJ��k�!�e���k%��W���y�`p���0�BvR��"�ʇk����O�������f���a���r;��x��ڝ¹1#2�k$rrڗv��x�潗>E*aa���FwΡ)�G@ ��5���ӧ��G\�K�3z��+�*�4({8	��$�T���ę��?�F�>�#����UDix����܊���fl&~[���FV?�C�;'mq��q�/!`3jeU<M���d�d�at�g����ԤϚ�X6P"<���/IcN��� ʞ�!��IU��;��u�ӂύ�`��2����$D@��uZ�6۞�^W� ` �7;+��v~3@����J��?Ë�᝖ɜ5�o(J��t=�w9�Thd�<�E��;C}���q%a�^��г����/�6�)��׎Z��&�l��pׁ!y����k֪{B����]xw�.�i�(^�"�9�������h�_T��kG�Wp��"�F�pV� �����1���^f�f%�-wYl��s`	�QK�
�1�	����Va���������\���.%,*`���!��dΈJ�fUc_(���@�7�-��>.XXy:�0����q�X<��Id������s����j���$�L�X4��*�2�v�C`��f%��Ԕ��+�]��o�}3�1�\al��.�ҍui�3�ų)i$��Ri��ȣ�K;�oy�;�)����+D��|q�pnm��E]h�/��/b;����BC� ����/m� ��Xa���+� ї��5�[򍱆�MA�.¢�hR��x�ߨv*i;�k�z�l����ޅ<1�@5���B�i,�5]�d���Jo�"[����z|q.y8�E<�Q�"�Υ��Y�l0�����]j	���6)P/��,$<!h[?B ���X ���]Dtם�9�$4z����	�|ϭ��[B��Vz�����AtG2���Sz�����lͶh��LFȷ'w��|�������m
���
����~;.�T������*��� n��iNCFB�0�)���^�@�5�ލ�8�a[>���g??C+3~ׁN���M����]!�kDg���E������?�f���5����_[�` f6jz��Gu�q�_|�u���|�20���UF�1RWd��!ޛ'�|�Lyk�s3�W̽�t��7�\���w;ļ�l��[&�,_�%QW���:%��S�`���6߁~q�M�A�VP%}�?d�Fy�RNfV��i$O7�O���lSƓM@�BTM������}��%�#A����;<������VE~z9�c�I��}�DW���mb�w��]��~��c�b��gu/�=P6\.�2X��a�8B���+H�Z��[��C�z�K5��=]���)5R�o"�����
y�O�WX�[����������zR�8��)Ys���"$irQMG���:�Wtr�X�z�_��f��(,N���i����MO�u�_�k��<1��e�t��s]��;9;���=���fCe�p��e8�"��`sx��N3���m,�( s�yq].��7���BD�?�xC`W$��!�p���������!�y,�T�uBL9ؤ�P#0��ψ;ț)�� ��ټ0�&���=��X�El"��0Es�38��L���a?�t@;�뼋s�$�z��Lmx���D����6sj6%�3ԁ����a�S�x�"@��業�~O����|S��1K{)L��z�&��6C
�(c}yDkِ���cv�H���\mM�*TC�����IR��4p��|�O)��@
/�>y�Tl+c��$7c�]Q8���`����ڤ����~3!t���\��9Ad���������K�5jĊ#�w�`���GQ�l�=~�~	�f��9y�5�|=h�m<7/V05��m�M'c!�F:�zL�2�x��/��}j���^��"��\+�u��,|,���?���̚7B��J�w��BY�v���c���v>TBw�3)��Ao�E�fM�%�r�Pz��An����>�Å��p�n��tqO�S����U�4���)�>��b�<v=��`�Qm�����҆�5|��W�Y߇O|��h+�+W�%���8B��T�]�M���������.�wJ�G
���Ef}b�zy|�A�c�sg�e_#��G䯗K?J}