XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1Z`nF��۲S�A�:��c4-���\�Ƚ�C�!�7<k���;�}�JN��Z�Чd���#�TAn�h!�.�O�S���L�"]CՋTB����U�����7�����_�����kʭD*u;�e�lɬ�c�"f���4qI��(��tPM[���!q�=w,�77`�>�)�]�g]�FA���lM9j ��8��ܧL�o�(��_�R"�V�(�� /kA��'w�8�����g�F�s�j��-F�üm�O�ywX�N�q���i�0�0�jgU��d ��C�,����޸e3䊚��:O��H����J�
k��X0��N e_�&%|�=L@�׼��:0� �?��t�>{Ǔ��pRYE�����u�+�]���x����e�Li�_)0w�D�^V 7��W�oƵ���a�d�9���KR�2wX�ғ���rx���<���WM��P]�|�	aP#��k5&�d6�Qtc�]�7�-s7���1���u��?'�%�H�pg�;�I�瘂��I��^�PSE1F-$'�'�ɴ�����RL�Wi䍽|���"T��=&��	:��ĒZ���=��B�/�P��5m� �{$�&��u�� 2�	� �z����h��0Ā||BF�ƽ2a�DgMUe�����jƼ2�ܶR ��=xf�I�bs��J�	�AǇ���N��e���,�"*tLظ����S-5)���bO���2�+��x/�y�k`�*��\���{�w�q�XlxVHYEB    8388    1740ŃF$e�>r͆54�L؉��c'��ֽ1W,m��qz�P�z�p�<cJ��vǲ������nR���w�%��`}��������x�K���n������\�ϊ_��EE�D�z�HM̂����ڝ#e+�G�=74ލ>Ƶ�&�zO��2'
���v�q��?�	�|fP���kC't��بD��;9À���{��5�2�e�)P�{��:��L};Œ�+_������}𲤧Mض�l��k����vt��Z+b$��Ndp�m�Q���K����u&�d���&�7�޵��)��q����Є���g����A����a_k�);d�I��4����	XB3��B��C4��CſM�l�D՛[�������8oi3�I�-f#��1�V��j}�a	[WG ��Q�������F͒�Mm�-�OK���A��[ȡY����߿�u�����3>��KkɈޠ_�ٸ���|Z1u�'��j�ʩh�����l�j����t/$�Y/�m<���H���|1�<���o\p�_"Ӡ��x�hLb���6oS�#i��N|s�wR뚞
2��1��`h'P��]�=gz�����H;J�U��5?
�o2s3��|����r�����t�Z�ܢ��9�FA�c7��с��}=�>�f��׸�U��4���f���"P�]P{It�ѧ��.��^��%�>6=?�^Nxh���WT��3IS��Ĥ��Dvp=r�{�􊤍M�t�=3�D`�O����&��}d�K���4}�t�3mB���KЁ���S�Oƚ-���P�A��̠���!�KF�Tq�Z��5n��g���q�4
$kqQ�����QV��b�Ă|�6�թ��;C�x�KU�E�esB+�/ڹ[��W�E�70���p���Q��G"�������赐(���.��!���j�/#�E��r��6K��gP�.N'4�U��'����p����N]�B=K�!ʯYh2G��s��\2h˓o.�5] �t���ڒK�0>�C��&��3��IMbkK��͒�|�d#)"!����No�ߡ�*�O�?��T~��.�����eԍ5�Nc�S��� !&kf?wd�w��"4O�=l�F8��4�đ���HC�{L,u��Fy^PX$�@A[�"�򎩣K�<1��7�G�^�+Y�h8��2kq� cSX�)jE|/=H�"��i�ǒ�I����3��n{ly�ԑN]I�Yz���7�I`
���:�|�$X��9�J������;/��>YaaD��\ A�i�KE(�	�Pl�a���(��D���xB�����'$]���]��*-`R*�ʿH�UYr؅���T��(��h�:(�I�Y>�^��GvRZ
�h#9z�,|@R��g�]t���� ����HZQ�s��lt��.���1���W�������_�$�PQ~β�myy�� ��A���(_��{�;'.�-�;�0��"P�h+M|-�
�aQ��>�1�Ur��6(�D�Z�6�[b'�hQ6S�]�m؈�X�wTj�*��l�p��<r⨴��s���l�IZLp'0����>۾��_��)J �Tv?�Ξ�X�~L)ީb:�n�|3�����v�x��6]��.�;[od�ٞ	�D�(*�o��t�h��М����C�h8��>���mdj���p�?D�!�Z���M�H�V��,ʼ���G�[���kB)s��[���s9���]���%�� f�ݛ72?��H�G�p�/������`�]s"�W�I�D�������:Vp����C�8��a^l�Λ
�I@i"�k5���2@��YP8��bj��$g�9�w)&?L�-�<�Gz#�9�飦��+%�/>�]�LzC�%~��<�`�{��>��QR��|�J�+�B��#R�l�2�L�̠\��8����f�J-�;��ڟp��	E����G�8��T��C7�s�Q��Q�����Z%�S���.�~���@!�HA�'c���P�ܽ+�By�Xz� (�B��i�MnE�&UN��#*�&�2��$��T�@7����|]0��HM �n��L0)�1OF�v@����.�^���;�h)ks�.�v���(�a��
};Q:��Rq��a�B �	/�PY&�7ߓQ�D�F�mA�����}����CǬ��|؉���h/�Io�'��Xg-Y��>~.�]���V�?$�8����Nb�?�R���|��hpA<��]���6�'�İ�0��z�m���w$Tԡ�/Pu��G=�92��BqD���7��s8`�Y�Z1����Y%���vJī;�э+�����9�1j�p5�u�ՙI�}�N:lߋ,i��cb�x�0��12���Qt{�)�������wS��Ň�����x�kc��@�$�E�~C�䙮^dFτ�I���,�i��aD~0$�դ�)ѻ�梥�����bD��d�#0f����9,t#���Q`��K����0h��;(�k)�2�X,� � ���"�ʆP��?D'�E�#�R����i)@�Q�1�y�-1ɤ�iž�r,VS������v(=�ևT\ꅁ�� Y�'T��`���!�4��\��m�c��'�z�[��@����{���UE�@�+7��](|S&ař���D��~�����Ǧ�E��%
�԰CC�ߎ���z�Q���7Ǆ�����z>��n�����L�4�d�GY�jB@�Ҩ-�YEUS0H��tV3G8/���������$V@�%�o���9�/dIzh�g��g��g�{��k�!D�z�e�L��"�l�gX�+���N�Ŝ��h�b��@��;藬��v��E/C|F6n�n��]�^�K�+�,�A^��M�-�zkoI��
P�ؔ'�q��"��d�P�$�akj�s�φkʢ�Z�.���7I�t�,�����]v�����t��K�g���rbZ��8&Z� `�Ӱ"�S��Q��X4��i��t,�i̓�1x�P�$�}��+���d��#?.�뾰B�3��	�BZ�%�����4���?k*j���o��U:	�]ov>��YoUF��[��2G���y��q~���S?��"	W.�����ʏ���}��h�T5�*�K&RJ�vP�����8�[��`�����'Ī3i�����'����Rp��2!�����`��M�|��/!��M	u�%�	n��Hώ������e�#�X��ۊB��C�d�,@����q�$5c�V�������6����;��P���8b���3gK�`zh���	��,`Sz*�5�?"+�޶S��X?4����-!K2���?���vq�X�u,���P���� �:�7�sWF���LA:b�-�[�tW�=�n�����x4O����WE�V�m�L&E]�m���5|$�5sŴN$�=��Lqp��(Md�	�Qc����
�`��d
�4���{*�um>g�Ey�6I� L�q���)��
?/���燔K�g��F��z��0	O��F)5)X?R+�9��5-�-����迕��SX�送�d�
 $�'+�큩�����5�H�T��x�Ss��K 6N"�@�m�����
y>H\֟�ΙW���W�`�?0����;��);�h?��\��!ݴi�@�̯"����TZh��ZIJ�r�\���4j�\	ρKddÐ&	%��R��z*�Q_���3����t�1'̨sǹH�����%�R�Q��)�����Xm�Ց�o�^Z�|��{�^q�.	��^�f�,�����l��Z�0�UW�
��������㥅��!s9�cǜ��v[�X]���@�{����LU�++	H�H���W6��2���#ϰj����i��<����U����7ۦ���n����R�����/~�a�G~w$Mw�J#`!����;:��*�r\+��69�W�Pw@@@�x.����aV�83�/-NBMh'�C�
��ݷ�������ި�n����>�
H4��qP����S�ڣ�Qi/+_X���j�ޒ��ʑ�uǾ�����b��*T#b�f4l��ۋ@qF��.F����s�5&{�?�b�5�sl�M��JޙR`p_�X⦦7*n*
!���0_��J�a�O����sH���l�qz�J��=Xl�!2���Lf�2i(EV|QH�Ҧ}țu(��9�{�0�;�r ��6!�i�O�ԙm}R���ѕ������w`г��M�s�Shú(	��G;_/Q�y}H_�u{Z�J8�o�JHlp����l��{9<$��� ^l�|gO�U�u���^G�F<0`Hxs�&�;��o9C�,
e��R������khS���Aі���0�Q�!��](��!��t���P�'���I*�����lث�lՎ�'�w҇6�<�q��n�d�}�3mZ5i�ew�,[���0ϟrusQ���-��hQ@x����wwz6�]�:�O?���-�#>���x�#Lf���[0��,*�)A�f�|%~~�˽���? ��l��j�U8����L���!�4�[ǪT�忠(y̝�8uzNV@J(�9ʡ9f8fgh.���[�iWe���J郇g����q8��#S�ٺ
��#��[r��Z�b-b@Z�JL���������[� �ҶOi�@�������Ǯ�.��
���7aŅC/��BX�k7��c���_ڊ��!��f�si��8x\�������r>OZ�t�PS�:��eN����:D'덮`+���9��6(2�+���/���G�-g-����;���`��tu���d1��u���w����p� �&
�)�H��N7���L5��5hN�����]^cƯ]���i�f%�Y�!�gǡ8sJ�@Y>#����5��qi8���P1�e*q4��=��#t�WEj]�zZ8Oڿ-˸�{1EEfC���b�VL)&.F}Gy���X~S䱞�un:Ќ���}���K=���<Y��`�%���"��sK������_����$[��Hk��o��<�yhH�,yS��:�Z5~�J���]a�w;E���������\=T�t��N
�K!���+lK�Ig�QnU�����g\�
ۧ�*��7$n�=�U�)¤)�^�ӏ�\n�oW7넅gęv7�p�E=��Ofn�6�#����&e���=��o�rPf
g���Q��g�GU@$�*z�e�0�VA����L]b4�5����_P�E������j���Y;�<ژ������>���Q��W��n
��>��ʎ�f���X��Po|�����*K��l�JkJ�[:�>@���-�Ap��u��M�QD_	��ٛ��v"����h�<�$Z�a*�&']�0�zv�w��a���Ȏ$�qc"<�r���r��l]~����Zo�_�~K��I=鈺D��Nz{�\�4��=n`K)\���f�@�e��:`j"�>��"I�G*��;xXL۩|L��v
�����<�]�|�:��Gzv'��n�dӈ�`<Z�@j{��9M�ݴ���R1�?�C:��*��y�b���dbk��W�z>}i��iaO`�'�E�hO�'5�x��/A�]u��l\Wő�,�:F�h��L��v�n����rn��5�{��7�kG�8�k�C_�R��;]^����Tpk��G�0�8��5��w��Y�V8,�;G��P��L�6�E?aϒ���qK� B���62���wG]�)��.��Le�0w��y3Pbv�҅$B�$V)�:E�G^��)9���ǈm`G�o�;	�V�4��uH_�p���a�1�o�B����[��W:�X0vw5��
!<�df�<�����}���Zg<���u�i!EN�5