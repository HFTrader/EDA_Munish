XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��C6��*\^�B�ч���0��"3�wF�&�PH'\0�VN�t6�;�}A�������
.� QӅ���c�D���z�6j{t�`��6��5��-�t3���p���A���^>����ڷW��5����7��Wilfcd�5���YP?�z�jR�ܻÒ�{�/�?� ��LG�a��r����$���|�i����斜v���H� 1�2n�D`�g)��rLy��wbJ�DH�@7�.��4��X��
 � �ЄO;�Ցzۓ�k�=�hfŮ��q���m�����N����V�P��F��|��'�!;��X3Օ?�Jи���g�%�R�}�M�)�����H\�5�6h�>R��a���˷�2����] /p�Dg�h|c���7調M�b��)eϮS�P���A*{���u^ؐ��Sc��M*�-���3�eN?k�#�B�`����`�:VW�L�ҫ�kA��E�e#(:!��K��=Z\����V_��_��$�~�j���(q珖���
J���>������xm���X��l�l�'����ԓx��"��[�zfK�r؇tlDtK��u��`H9�>���H�MM�u�'��.Cr�kB���w#oHH���rӧ�\�nug!�Qqz
0�a/OA}�y��������Y������s�N�L�1�x��P�mA+V6��e� 喢l�-����CsG#7����@��'C���1K^v+��,�k��}����;rG7��v;9��XlxVHYEB    20bd     a50��p�^C�+W;Kj�qw+{�^4�RVn�Ǎ熁W,L�m���Y��u�@�T���:}�o���Ian#�f�JR�v�9}�G^��K�Z1�/`�IґC�+��5``3�X��Kϊ�	�O}1���Ɵ"��8� Vu�`� �x��h	��a_Q�s��֎�P<fç�A�=y�w�h��/���k@>�}h���������y]0�9�0�9YjLo>r�(�x��M�$%/u� ��J�^p63T����yPP��1y��@�zZBb����5^�W��1���5W���11�#9T#-�\GyX��~��u�ÀvF�`
�5	zA���"K|�K��*�#��.��E�L�7���Wr��;G��N��+��p��ؠUX�ŏ�Kq�`}J���+�2����=�B�=8�N&������@q��ה�IAmP<|6�U���Β�{��#�,�G��K+���\r�(��i�ڃ��*���H�HJ#]f����FU`�Som�kFf���QO���)�� ���vN}�I��^�"�{�b���B�4�����h�7�;�J���:R�����.J�������n�~)�uo�F�[������`�Cek�\�+f�f�-�&���5��;�ɭU+�L�/�h7��%*^�/&�n����Z���(\D�Nׄ����Z~F#4�v/Z1_5��1��3�����PJ�d[�
ꬅKЮ,?�{��!�=��N�vG�!r��*jf�@��9q����a2���g� ���-���}ZmV��u���R�pZO+I:j����{�����a�Ղ�
�˷�m������#�꺃>^l�LT75��"��>cy�\!�)��� gqѥ_����mCU�]�&m��dA�������F�Z
�(p��;Ϲ*1�[}�;�7�֥������mf*j^?���������|�s|p��ڂ�!�si���̠�˸7;x�G��$�_�T#&3"BN|�� ]_�?�u�vԍ5O`���K��G9#\n��"t��&��iCq�IcӃ�*�p�������l�0�k�3�F�G� @EVN>�?�ᚘ�מjl���:-~L.�
�����g ���0L���~��Uu�|��dzC�ҟ���b������|?�R�ِ)�*��A�qGr�����BöwL
Xs���z�uI�j6�՚��m���4Kv�8�_�6=oWk>l>K�F���$\�"oe�P����蒟���@���m�ol�
{��%̠ǅ���3EDW�<����ט�@��qG��B5�I�wu�B�qk�B6�f�Nl�J���}�;��o���tH(��R��Rw�)�GS���B��+ ������85�����7���j��OjV���� h�_�L�3�<�*bO\!�-~q�4��an�
,P���x�e����ϴ����z��8�(M!���e�(+z���%�,�17�t���h\��'i�j�wǢ�-*��/m���.�.d9��t����+j��k���ֿ�t��筚�J7�����:�د|
7��=�M8B�e��6V~�9L>]�����n}����Ď�\>����g+m֬2ڱgKi,乤���u�r�6i���%0��߶�~j�h�N�b�G�6ׇl�.�dV��v�_�8�ӡ�o���(�^�� *	�PR������rKD���|."� �Q��4���p��*qU	�D��!8��Q*s���l��r���+��0�`!���$��b��W�φe�#c
�L����s*���z���"�����k[�i�M�jX��i'0��G �Ec_���S�L-rY�Gm�$����I�e���D���!����`�
VAu��p���ff�N2uT$ԩ��inFT��YRn ��X"w-9M�MHh�����?���ST�5!��bvچ�N��V�D��_���r�Hb�M�A%���jn�԰�1ƽO�VأOO~*�|�Q@�`m/e#�u?6����`ऊ��ط��!{~'P5{�\B�����,}?��t"��H�Ѣ�^�*QB���Ye�S;K�0K_�<�C�;����kN:5l���Ъ!Og<D���d��|�{��0�j^�hJ.r��^	��D2�hH�m�NU�z.SK ��ʙ��:�~�&����&锟�Q����'����"����o��F�$
2����N��P����r؋��7��p&J���KM^B�%������;/,�"3��.Jn$�e�IG#���P�*�&Y�hhș2m��l2�æ�q\H�z	�ӰP�hi4�H�B�`��U��Q #)��ＣE*���������l�tFK�uq�M�'_gB�%�oף�#��N���J �1���|ϧ�>n3�b�q2��Vf�x�����aCX�̳̊�Df,n�Y:e�1#-�JSq�)�h�QI�����"���,+/`н���'����T���n��*\��^���-UI��c�7��L�_��Ds��x�^���/������y�XS)l��<����n:-i-�9�H����J�/P��@�j�Pa3B�֐�