XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��,�W
���3֥�4X�h�hJ��`�����Wt�}
.�H��������J-�.wc(���}Y�������.�[/֎�M	��v큹cf?��B½�Xy l��I��h��e�����o���D���ɢ����Q=Zo1����]DB���Iq}���<��^ڀ���".�	L���~��a�����'Y�_�od6�\����3�1uj�,Z{?����r��}g�Q�!ͻt��_�/�yS#H�3����O��]lV��m����I$d�3}��S% �v�V��s.�dѤ�-����RHl����l� Ǹ��ó;��KMX�.:/���� ��QQʿ��C�U�!��'��R� �4hl�~�#߰Ջ�X�ܑ���#&�ɏR>�����ӆ�!�O`���(�@�42��ۏȽ�u�|�n���D��fx��G�حy�������5�=E%ӄ0���}�ke�O�*?^ZB�\�ۥ��OdTk-��ȼd>e�l<�$���2�?����p�)�YM���T�6��ե&l8�3�!�NUp��x�&����p�ޚ�Q������7�}�颰8����P����,��lL�7�Sf}WL��h��{4n�L���p�w��ӧNP�c�������<� ���>^��hʣt�_��?R8))���f�F)ֱ��8��[�Aޠw����B(��OB ZôD�+���S��!��9�8n��X�Uő�����źt�+�� �ÿ��{a9������l��T�XlxVHYEB    6014    1840����Is��Z��h\[��2�����ʞ_��� �7�M�>Ә�K ����[}͔4e�	�@�P�P��9�$�Hka����Mh$_����'�n��x��D��&���]h"A �L�La��
��*'�,"�%hw�[nI�v^9!�fZ7eP`�ɶ���iR�3�ˆ)U���=Q���ּ,�SK@c@�%������v�6��uvѻt�t;N�+��p3aҟ!{�!�Z?��8�D�����|�	�hU�b��j��Ɓv=� \~��$�<v��z[>�py޲,��IS�A��\�!�H�4�_2yj]����1-�U�TG�
�٧B�	�u�YY��X����+�'����MR5�9̼qf�ø=�F���
h�,<X��T�bidGtU�e� ]��$"�,$�?<�fB?��׾��Ǵ����&�(���-�,9j�+�c�Њ�ϯJ����O��B�X�x�h-�4xndV�耷Fx���'q$+�ĉWƖ��]I4N�?��e-���� 3%���ʙq͓�k`�m{��+oy�[��C�1����T�qkJwv�Z�B�+��O0�����lv��S�D�tT���@nCt��s���1F�e��c(�!����pu�``�h�R�P,�ͪ��!���"-d$ԥ��#���'>��nh�n��뒂:v�'J��5�q�̑��p��d�a�9z]{(L�0�cT˔�`��NH-���?��g�'8��əf�c*��U�S@�/A3��%uF)&�k#��[��F�Ԃ�@��]L��R]�U�#��~m�W�ɾ�Ә��o���a_��4��95A�,|UĘ�u�a�<�ьaL�R���(p����Y����z+m����s�۹'�F_Ѽq�RO}�M2Ҽy��4 >�h�c�{]��W�=�Z�R���c�>�N-�>������|4'$��������(@l?)����	#�p�;��FC���e��[�v�w�H�^O��/������e� �Ӡ
?��	]�9I5{�g$%��b��5S,�y�������O���+�����?2fW���&43�T"�Ӽ�V����{�]��p�Q�$�8��:�rv��R&���{0R���;=J�k�u�Z�a�$����=(��K�GZtc�X<�0s{���y�7�@���Q�Cx��o=��?�et��Q='�,ȺA&o�4m�1�����D2t�7�+	�1�//�{D72���W��U�&l"}|��ܜ	��n��6-iQ;WB*5����/��>ǳ��" ������-�VV�i���M	lY��\,ohѫ��8
@��9����[�Q��^��2��c@���%��Ki`nA,#FS�(e���c��)9��9�e���{��;wa���"<�v�x/p][8������o��2��K/����
���埙�G� �;勎�,�#/=,�6tp�����4�i�'hj����0���E�B�!gGh�e����]��eo��������N�^)����"Z1(�k�H�o(c˩%�l�I�Æ� ��P,���@<^?�6�ڒU4+ �;�_]���e$�����-am?}���$�ڷ���۾��d ��z�`Or�_M]� �ؔ_�ʾ�fk<YRXc�Ϊ��B0������%�����X�������XG���ǟ���~AP��2F� B���v
~���k��9��$�bˎ��9��?����N d@��<)���#�U�3�%{����L���mрQ� �+��v�6�aņv��MJ��ϫQ���q+�i�晫7�n�
aB*�&\�O�AԂ<�9�""�#��0���-hD�����^|�g�o�$����̣g�8����䲩�#,���:�����U�)�p�ί
91���K����\�8p�0����o?����*.�i.�u��be鬛����?k�c������ -b��{e8�1f+{sLĠn�AU��!3���-h���7���V��s;���"������!S��u[]j'@T����=k$�\�;q�G�2<6�x�|���<#��R'�5J�>,�)Θ}ø�dr�4)lU<�tM���<�C�a��9�4��z��� ud�4�}K��辙[�^�|�0sѮ�]}���ʝ)	��p	�
4�jO�'���@@�S1h&o��_��߬#E��p��v�%�T�)���eZ2�]�,�C>������jv|!h+L�f"��S5�V��D�.��<w7�����hI�' ���Y.��D��K���2TI�m ��cS^�X�O��Y�V�,�lP5ȿ��_�tU[%���H|$��G�.����ᥔ��8��j�G'�1D�_(��hO���6�G�K�C�7�[�� t�6�,n�Y���Ž#���[��22�7�/�h��;����Po��}ȅ>��;k!�)�a�b
!�g6�6�2t�a�Yl����un_�B�@ـ��'�T� �#0�q��1ʓ��1 )����G��uPm4�s^_�|��yw)�4���S�Q��%������)�M�4�ӈ�Hrs{�Gy�m&6�2R������T^قDs�7z&W������7G�KI�k����v�o/ABj��*j��҆	��

y&�<1��zm&�ւ0��/��<�&��1#H�.i	oN;B�*:2VD���b�#�(�I��$&��3#�A�}���0�����,�+�OO�@��9�X�[OwE����,y�sXΰFY��,�����p�t0�F���_��f���&��GHPܬ����eI��(��:����U����4i��s�������ĳ�+��E��r<Z��K�dn?@Ԧ4ښ�l�X+�S�`1���b)ަ�a7�a��8~���;����.$+�j/[3�0��8¯�z���d�5�A
���z?�F�D�����)Im5F���t���iV'=l����)��d��J_��i�d׆�5A��[��~�%M@?�*򖿞��)�u� �Vv�:��UI��4~�[p�39��CY�$�ul9�2�¼�3z��{pP�$��5/o���x�ǳ�S����{���܀f����ҖX}2��ğ;��U��F;�o�����wGưb��6~Qҧ�
��6� �Eu�F�)�%��tx�k��JA���[�N8�l�W�O���H�u�m����w�0#�<7fQMb}7��_C}�Q��� 
�{6�/�5X;��Nգ13��X�f͞Y��'z�]�妉��O��V��A/ v�����8J>D��mg�ybY<�>�c90HҠVQ�؆~dIB8H�(~ C��&����g�U�^_lD*hD���aNG�d�IF�� � �	*��MՉ{��G�D��]��"p2��C\�G�7k'i�V�'�.����s���z�(C�ō$�Y>:�;2�L���\��CӉ-CӲ��x�[�c}D��PqpN����bt|KO~U)~_�W�Q��������in�a6ԫP8*p�Ft$�vߜ�|T/�d������x�E:���`�)T���)C��5�'���N�8�s[e���F7M���|F)��ʷQͥ���s�SC���{�������Eh�|:"���FG��*�LN����{�9ۮj�]Qc��܏��������#+�B޴��3��7-,C�	ٍ��C���ud��oq�U�Rfq?62e�)��t͎�-$P�wT�,��LU�~�?�� �������(j�R&^I�c�e7�����W�Y�h�7�b����rS� R+����g�ؑh9Z�5��� �~Ì&ì)�쯖c�z���y������򱃋)v��&1��-�Jۜ�"����6�HJ�屘S:��3o������S�v4�*
 ;=�h.	^e!^�BMv���q\,��5���MW�x�lzC�x������\o]�V̥G(����`c7��)��2,�$&[�zy���O�ݞ�Iв�#�4J���@�C�H1���M����5cP�NA�r��^6El(���3_�K�%�����~5N�L������0���&��
�+�<樬И��A6n1�c|x�5n��V����[p�>�
����ǲ���Pi����ܺ�l�5��G�@�����m�e5��v���b$xm�����#$������)�h�X�B!0�Ag[PX^,���n>b��`�����V���UjZK�
S?����KH$1D#�S!�$m��=莩{� <�@�$��}��섎�H����]Ӽ�`�\���7YN$��@X�\4��{R�g28jٲM/�7��f��Z�`�j�K�xT�>�uV��P���(8P�T�{�b;_�(��5�g^�Q�`@tK������&<�f���"��E��# �z;���UĚa::"�;���g�ƒ������s�!�dr�����
W`-lP?�ir9@���Z�U���{@�� ��ʣ��mh����gk�����v���YDw=��oy_3$��.���\ϖ[�kh.�3�|�޾1�)����^Ȍ#���K@�;2,�����Ŧ0��*ҡ�Or5g���"ኍǪ�d��I�.jp����'yԤ:��y �K�j�;���k|�v�'�W1�f�PL�A0.1�ڛ9*�!DO�u�_�F����Q�-����R1Oԋ��Ì�
 �#&���`ņB���V��#�YZ| ձ�N	���
�:ܧ��te7�ҽ�
�FVl�	���]�y�b��`���gf�aX��<�ۨ���P<_6�q��	 �Y���Ӝnk�g��Ɉ����8��Wy��էO��%-��l>���o����l;ײޓ�aj
�ɴu����-�q�#������j�;�z��w��ѡ�zQj�)�`x����x���1o�ShO鋢a�.�!j�ʎC�C%����8�����m1�1e�^��	�!�=K���c-A#��`�m
��nk�!+�E�L����o�U�^!^���Z)co}xqx��ס�>�U�,g����YfӾ.�$X?�p�-�n�y�i2I�{8kfQz�Sᑖ}w�Y+bӸ=�sk.u�M��u�K�3�?���2�l8��#2��=M��֕w;���8��۸�r̸1�k�Ŋ�
xem���W��ry�h�����teX��$(ayu$.���u]�ۿ���$A�@�=~p��|��f�z�~"��^��'�]��6w�Z�*�N!x����;����I����z�E�].�bCD�Ec�ɉ$w��Y�j#p�)�s��w�&��Ԡk����,!�t�Q�d�@y������-O��[�����	�3�_Ϯn�NQ�{@�I$rUY�Z�I	Z��m�����A�G�@v������nQGX~!�{f!Ɠ����[���}�t���E�|7�ڞ�x�y�?P�����'W�b8�Pq�{��9�Ԧ3�o��K��4�bO�E��y�ϭp�3Ѷ`��Gv Z��ґE��������[�'y�K;�u�ĆqGς;=�u.<rE�f������Hn6���/�K�=��?>;�	\}�Wv@$�a�b�Ӌ�q���t�,��o��o�l�끅�)~3֝�,�8\y���G��]�������?]����ќ��|�R�O��n�0V7v�V��"�&I�"!^����L�ZfS�;~8��{�b�lr�h���U�iM�\��G.SUL����O�tI�8��!iZL-�=��+I����Yxm��8�9"b'����'���Q>�U���j�����-)�O}2���֝��W&l�6I�~c�ǯW5����&�Y�6�#w��g�ų������ꪑ*��(��ҝ��V�MHV(� Ȯ4��Hk�loޟ�:q:��V�\D���M�d=� n��f���DVdAmg�X�R�慀�"��Roɴ�S�W�Hu�i�b���.8�5`���Μ�`6z�ӊ"�٣Rc�*^�\>e[����o���s`�5���U�+�;&4.�0�b[hiN/H��J`�F[���#�w=.B҇&���]e��:���aO��t<s���wDl�'��έg2&{(�ݸoЌOd�B�!Tn�E4Ԝ)����p�C�