XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`j+��I*겓W[�B}��ѿy6EZ߄=P>��m�cy�-�ȉ_>�,bʹa�g�Ekz����)nc����
�$�o��.�ex�O�=�C���qx�1�L#K���q��ķ�E՟�{ʠ��/�^>0:b`�<�ÀB�U���v�4Y���\{Y̥h��f���G���Q�O��v6+⃵Ź'�Nd��֍R�{����LI�%��]H��W��x�f��U`�i���$<PX�A�3�O7��)��4w%��.k ^Eb���)&��a��,eŤ#w����#�b����ʀ��֙LC���!��[�pr�a_	�H��I�,�^^M��6 ��S_��u�Q��?��k�BGit3l�.��@��Jy��Ex#@�cS�D���;�
�~܀B:���%����E�j^��Z:��q��bz��o?9y��)�ݕ��\>Ώ��s��X)y�y�$i�J}���&�]�f>�g�=|�{2����)�[Ω�-l��۫��/�o��(%��D%��y�uy��aC������m�d�>89��㸨�bR��2rH�x ]�.UdsG��{J�p.��W�������������=��٦��8K)<�P'�~��WՀ}�GX��%|%�۪�n7h0���n�)���OGs���t�X�$��9Gה]�*��l��w�i���K����9�l��n��1���~�� \#�V�\�@���'�7Rd�T�����N՟S��WwQ��$��hmi�RX�6�VXlxVHYEB    117a     710��?ɠhڗf�w^�hh��8 ��й��p$d�Oa���%��+E�#����K�֍�iQX�0�C���D�x賐^��Z�m�= ���(\��,8uBdYb����$~[�mhG�M�
��1#c�1�j�< �#z�麢���~E����,�v����D�XrSg9�����pYW��h�F70�����g�%�͐���˫�Ի�t�Uq2S��d��8/KyEZ�mV�z����g��E��T,�	�Al
��&��ΣcX/]W�gO�(R;hR���hc��j��{B�1� ���iL�$�`��
]�K���3S�ڢ�d!�X�g�~��y�
TT|d�;YcKW(�a���j�t֡����։�mxY"L�d�(�%��U�򩛇�xLUEf��RE4��P�Vz�b�H� l�s��,.i�[���^?ְ��JhA#Oh�����<�' Iu�p ��~��S�:k����Nf#�P�*�mDL��s@�Zu�N�s�/��w4YJ.�X1o@��z};3��ط��N(,1�@(:�	2��_�o5.�n���0����\���Sm�g ��p��s0��Ћ$l�����y*P���R�Y~R��E�xk"��Nd�O��0d�V+�j4�\�h_�oB8x��Q���7Z����A_l9�$tC-�i��%ޛUN!&� \�_Wf
�oG���'�o&l�QPq�n��Q,�4ZO�x��V�����k��-_s�i����i�ήx�/�H����_�3E1�6�����ks��]��ظQ��%a��F�h�7����<hZ[�y�G�͊XG��3�i�i-W�(<��s��N)��Zs+��G�%�ek����b��n/�F���G���F�Wd�ω��t�*��J�g���L�y����ڄQ(�e�*��h#��]�fpLw�C���m�C�~l){��AF.!O�}����0u��ȭS�SJ�*�U�����F��(1G�)�wum��i1�=��5�GC�Ctx(A6B�j��zr2���w�߭���b�����6�ϺX�Ў$�M���S��?��eAC�����;�i�3���T^hy̥ (6�ry�h2=�XR�e���6�����rI尳��\V�앒Ƴ������I����=��q5�p��JsB�����w���/�I�ܶq�� y7�4�l�)�+��Y/�v}jU�~<����j�/~%pCk_�J��s�޽��r��sDhۗ%�m�$Y�^��n#�0媥�^@��+�XFL��'��
���U���� r/�hh8����{K��09Zr1���S`�+	�ji�cg����lK`c��{鸱ݭ;��j�p�t����5�� Sˌm,G�3�pw|TD޵�!�`^���U:��ѭt/����i�W+Z�y�V�b6�~c)�ܯ3��F?Q��F�����p����=}%��&��K<ƈU��>�&0��ˇ�Qg�4�2d���Qm��+�s�2�o(��j���;��uK�=��lY�2�bE����K}�x�U�@�>�8�刮����e��"�gcc�<M��s�&'�&���ɰ5KHg�D#ݛg��Ĺ��Y�T2�Z�wN姈~W�/���ޯ]��S]΅w�������h ��Д|�o0�ϐcW~�+��o����/h|��l5�Z醖��,����<�����L!�����I���!ۭ�< �B���[kj�S�6ԟq*�'�ZJ6#��l�9Z�2�Q|Ȭ�.� ,� �vu�s�q�[�