XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��]6�]�g����Ï�4S�`�$V/�2 ȠpX��u%Dz|��:�E���爧�@ѹ��⚻>lF��P%v��&5��j�Zis'yқ��s�r~_���i0��穃(7Wі�>O���>%,����7@���2�[he]
XuX���Zq̕M"�E!�.@�����e56�Ej����*������ļ��I3��j�:�Qc���5
.�!P�h�5G�>�>ʩB=]�7`��i@�D��(��S�R�u`D�D�2"���r�g%<\<�.��Ӥu����e���N�Z��Ì=HK��:̥�"�3aE·�����̿��b^�g\.��S�J	�7��TУ���G���l����R�R$m�_��'�a��À�i���pEf�M�Gx����)��dN��l��,p�'�ThH��"X�d�� �R�v�z���o�<Q_7� �����j��`����0���V/m@��(u��Y�iPT����㚶�G�I�-�d�#|��%��J��a��i�q>b
.3��>��+��s(�k�\E�˿Jf�������\E���S�� ��u!2�9���%҃+�S=��r��g����g?�Ӭ�d"��|;gY��.%���z�7ȳ���]W�C�\�q%ݪ
[7L���D��Ȱ���}�
�C����A�jA�zE�Z%g=�zhۙ�/��8��@H{��V<a�/�ոd�|L��
�L�xꛜ��vM����_hR�獱6~]� �^)nr3���XlxVHYEB    70a6     b90��L�rK9�D� �/�O��J��`i�H���19� 
OW�~q8�sِð� �<e�ZX�l+�lZ��B.W)�#������_6����D�M��c���D?��O�$�!O�lk�3cx�G���ȩT��Pẗ́!����H��5|�L��s�
�@"ݷ�I~�5~ېҹ�s�x�B�$�����2h��T��w�c�01��c1ڔ�������Ѫ���e� ^����q8�s6N_&�씌���=�Ԗ�ZK���3�������rT߅�����Y�-9HlU����?���C�x�:��ㄇ#s]��X�C*�Y>�#�Ex����Et�.����;ǃ���Z����?������*���"��z"kw1���rd��Z���{��F�
F���2vE"���YJ��6O�A��#�xI�(�ḙ�m�Ŀ������N��F�莶���E
!�~�`�2�bJ��rf�����j!�����5�E
]�7��U�۶����w�]B؈W�!HSV�)F�-��\�T�0�*�GE�(�r��S?R��Ċ���-�,V��3vS�l������8����d]��������д"�Fn��Af��>���ad�g��vr��qyfL����E�Gb)4˓��t�T5�u���z&�⣡~��d2�}uA�J#X�1j~�.}������E� �]���p�v��Q8�B�@�՚Z�k�/�N���V6<DH��͆��H�%��M��x�b���:�|&)U���:q�`ly���8LN^E3�=��W�)� ޑH!y8#�y����5�K9����NY��u�&���#��{Z|�@� 9H��L�ǰ��k��Q�҂z8�X��f�@�z~�i"�@A.�c V��5H~�҆h�h�˿_�-Rd���j��o+w�һ�L�Y���ˣؑ!�"94��>��*o�pQo&�,�D�L��T�-����/���b@���dh�1A�l�(А�g-t&�3�z/��^�̓Rw��R�i7�Y��fj��Ѿ��6ε
شZ�0�7�G h�,yl|���-\.�Ϋ.K	�A�?U���f���k��O3z�/�d"+�z/�wI�z�����l�e'�Q]Di�~6ҋ�l�8x��)�)����@&�0g.n��\�~�!o����Jqb��;�q& ��[1��7�3�_��l�%,��~���M"��w���H�m%����I��&� .�^~?y�g�.�F��ɺ'�K�T	���u��� 5�=D�5]��.'a�P.�L�.c�Pm�<a���4F>�<5�������A��P5N����!��dd�U㽤I��ͩh�D@�_x�PjUD6����	O�@w�����q3.�~�fS��|�ܞt�Uq.20��(��}̈Ղ�����6��sI/��|��洛�́�;���;q�jlݖ,o�C���y��6��.H`Dc��kf��R=<�����Z`S9�����ݍL����\;V�-&�Bv PUem�+��i&L������u�|Y:?�A�H�s�}��sÄ��}H��W�`wy�������/L�����$�+a�z��c�Z� 1��<M'h��h"M1�U?����1j�2 w�>�]��%�:{1q�bG�1�+����Y3uD��>���cQ~��X?����o��hlDf�`Sܚ����fn��l��Y.����V�j�#��T�Z,�Um7��'Y�M�����#�7�_��TO��-�{/Q�u�cP��%�-�t�78�$ɾ�ƚ�jP��pn�!y�� �Y�q���Leoj���o��"���7�1�C{j$7g @�k:��ROO������Ȟ��4f�8���w5I�/(J�@�3<�e�&�T&�1iKu1�b�ǐ������Ls��>kۦ�.z�K�N�w�0��4`��H#T;����W�BFTwHxU=[`W�� ��M�1���o$��_��6�k�,/RĆ�����f�x�/���M�us%�-V+�Q	�o�V3P,�F�#'����U�w[��K�^�F�`��Z��.PE��R ���.�]ў}Ayl���!){��<=nR���VD^��C��TKoQ�t��j_�)��%ԛ��rr&�Ζ�$�9ר�O�:3��dL����Eq2�eD'�l���Lr<��R�C_���F���IJ��b&�`~�ZLl�����c�f�>�F�Pi|@X��ޅZ'q�ٚ��H�ْ���#��XWƪ::�}�J���9P0	^��*cY3��-����Y��������d�cR����:�eUh�w(����\s� A���碜��1�Hg�ys��4�1����v�E�+!,Hk�o:I��a��jh9UM~���8��R��� #��pI�Ó>;���q'/���+�!�\�fv�r<����	@���#d��|Y㎓�;�]x��k݂�8�b�`'@�ٴ�R5��ѷdg�:A,Q�z�_�O^`�Na���&��Al�յ�cd{BUCp9C>\�W�F�퉶���x�a�L�R�@v������I	���)���9-B��˷/bs�җ�i���z1	,��2���MU� ��6֓��J�΄�d���)	�@T�̤N\}�.����wAF�M2�C)V@�ȁo��˱*��l�l�

���V��<(L�� ��#�A����,�����(���RtN����A�5��~i#ah�{k�������w]D�����/G6}f��H�����↊����ugk	B�E�q���?&�v�:�;&o:��	�<��i�b�3���UgQ5O��:q�\�
�s�Ke����:E�cji.ADa�?�L]Z/0C6o�6���W^0`bKJ���e_���V.wԍ�>�:��iV�x����JQ����=O�Xs�� i�P�
���