XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ٔ�=i�*�����!�8_SXM���ĝ_��=��f�%�������f��ʽ~�4�v	Y�7���=ޫ��J_�O�z`}���,1Vo�9D��q��6)�gT� 	����qBiC��`�a}�J��!�Dɛ�UX���N�k!յ5��i�1���0��C�sZ���Nӽb��� 
��Y����ʍ��{�9�g�f]Xnާ�Ɏʩ��;s��Z�q�h=�%&��TSgB��Ab�4;&���Y�r<��wqG�@�tE���sxJ���o�A��JYh<���%���i0�mq�M�6��4$7ޒ:^��M��H5:�MW�#^����Z�{*}��Kx)M&�������E�(��X��nF?p�k����N/|��Ι��7��W�����b�bc"�r�	�a��H��א�>�t����L���x�~���J�³��M9pT%�;�$�ڿ�3����ŉ�h�͎�|�:w� Ʌ�d%��q�w�d�q"'�C!���eN�XӔk���rff��"�{�
x�f�������"N�@���M9L�p.�Z�{*@�O���D2~1�R�``����P���{��2�KV6^�ʭ��U�+�ALp�
�gO������)�C�)6���;|�,En[����`��\��b���=!����?�M˖E��k�e ���pʫ�xy��-I|�����e;Qˮy�{�ښ~��Z�,�Q�a��@������7����%<&�̤���`3iL��c��cF0��WXlxVHYEB    a037    1fe0ˌ�S�����x$q�͕�iŏd�a@=�'��f��_7`,��������|6Zj-R�\�Ѯ@��w�'�\��?2�f��i05[{����\��b��D�N�k+�!�N��B!6b
N�?#��;���A(e���]�CS�n�B3!��4=��I�.��ܷ.��zOf�����VK��Q��u |߂f3ҫbW���J������@L�u�A$�%��p#!���'Mܸ�8t�Ed�3U_zn������F��w�Ik�c�z�$���:0�#�ؐ���3E����q������DC�B�ڈr��X1�F���+>���"Nu�����k���3q*n����ӕ%}��L����F�"�O�����s#ů�J��m��f&�9�m��׵�HZ��|P�Dyѵ7�}xJB4lV� �p����L�K�W�Z90�!��, ��_�rz̼�ZL<S���P�R�%�v��a��{��|E1[�ǭ}s�)���,��'뜶w��8�b�M�R�ݻ�
�N*�0]�H����kѠQ�sk�\�F��;�8�4f��"�:#̤�?�m�G�6��j1rMv�\�[|dE]�b�.0�bkItw^�$�)�5O�P�o.�|e�0���Y�O�b��J���Mjq�n��W����/n5����Ul�9+�q�ë�)?�G}я����iT��F���X��e��>B�m������t�IW7�f���_�[�(P�Ւ�<��t���3 ]�(��B��FT��$�q���m��Y���8u�"O�c�u�=�m�� 2�t��#̂',�xEW��&�m"~0[�#m#h�:^����64Nnq��n.D���V��ʶ��w��l�	�{���I��L%� L��5ه��P.�0��S�Z/����#0㝹����#39���雲�^/�v��ݒ�ڡ$h���|̴���o�8���ل��fn܌�f�^'���|�f���3��P�k�B!J`�\��ecp��#*|q�oX����{�&*w�{7���5���\ց�<����6w��a�sqct�,HP.Ji���T_���;̷L=ͪ
���(/���£�� �q�uZ��`�B���Hi�@Kݜ�	�{;��
���.<@+$��J��0ׁ��mS�.��_0���}��P��BtgY')X�m�V�c���9��^��x��D��{�}7+' (bC�T�1�����@�?1��_0�Y2sB@Y����ޜy��A�*Gq�:~3�t���q��H�m+4])��$��,�w�1"mv��,�ΐo�K�}Η�2����:�g�9^�w����?��-uO�nFgUi%��
Mz)_�X^7�UhYC�{�k�M�HX�YzD�A8U#��+�t�\ĤS��k7Ӝ0l�W���%|ng�0�Bk�#�i���`hN0������W�����C���!_e�6䎵����p����A#:��}������/r��v~G�&�cGV�$nE5t�u���U��^���h_�$���5�:�TfY�Wꂦ�?���⡹�P�K�L���Q<7rt�/��N<��"���W�|�4Xjye�ݽ�k��e�P�B�4�T>�ѰU���^Hx-�X�iO�Ԯ*�����X�K�Ǉ�JM>�$�0��⼈�n'tmҺ�ĉ*P�{Oβ!p��Ŧe֎h_��MIl�f�|���8\R�w6���>y�`�1�#�fN�a�@�EB \���_3h��k9�f6+�X*�.L�#�m��0�t�O�ɧ��{Z�ٚ/����⣵�k��ewF�B;Ξtbn�9)�ade�<q�z��9�Y8[����fߙ�[Z7gt^Ԑ�׏gNq�Ra�-ڕ>�c�g�/D#(��\���;���=����xq!q�t�$&��CO:9Q��j�8c�AԚA�~N��N��k=�l�|l"6-a���01w���H�)?s�+{�%�qx�E:�Nٯ���U�l�w4Q�RF�Q�������R+��G}�_���\a!�(��żį�qI�V۲�;��stk��//C���D?��F�n_
]���'b~�Va�D-�B�e�ON�*@&�hwT��
���#[��+��������/�oR�R+�l-3)l�<���P�G�9B�8z	�3.���H�������z(� oq���'���R�Y'h,�~�2Wp9	�Qm5V�����M
��%r��.��!)�(���z��x�%E��i�0b����Q�uS���B�f���D� �Nk-�%#=0/�E�{���'x�ٷPr jւ����!�q(�l2h��~Xeؕ�^-Y�n�:,����W�����9�8�!g�����#�%��
N8�&D��&5B D���q̉h�7gEx��ɦ���p�mj�m����%��h�b[�V�4ѿ��k`��Whg�o�E�̊�=����5���`&s�O�m։^TN�\�OB��R]��|����밵7֨����3��'��Ю}�w��L ���ef�F濳�Qk�=D{!�{2l<s ��u�T�%� �����K�t�`,(؁������CIu�74��nZ�8
$���36��iX��f������!�?��n|�fq.O�r_GW��B�f����`��_9=��#S���� 	��^�U�<�=�%FJ�Ұ2�n\-�5=��������OhS����l�Z�Ug��z��WU���o$zk���2��e���4�_��.HܤO�����+��[PѰW*1�Q=��(���6�S�A%ѯe�N�Urjm|�KQ�bؑ\�q�Q��t-���k�|OPQ_�]#��hȃ��>㱎��ۏ�������]�[\&y6@5`���[��zQ����SõW�����v{T��<�Գ�q�׻o�?0�D�"���9�^�iRO�B"e{�כx�5f�թ�����@���հ���<��(��$,J0WO��ϰ�6�6��c��S�Y����͈��a�$����,��4Ib��@�T����f�E0Dbh;�|��y.sKa�"��B�sĤk�L��âp}wzn�0FhX��
��R��T"�����iS�^�F�w��Z�ى�Ը��[�!�� �]�ę�N�4nFF��j�]�{���V�hə�0z���-[�J��lp���򴰲!�<O��	@h��Ղ.jn2��!�@�Qb��:C�(vb�|�� +�o�g��N�Igc�W�$��!�5�ȋ�W��V�9����Fo-�0�ڻ�oދ�Jl�"��:�#u�����;�(���?c�Ko��S8���３Eg�8�^W𱗳���Ǩv����l�v$�{]�E�αn�)�У}6���X=<'ΎN�S�t��5M�;��r-�`̦�|�wf��!�f��4������g���U�ZL���UL^��XFA�ʮ�QV�%�����Ҫ1��x���tC��ك��_Bfk�)p��a��0߄�y�'0G�+$#�h���[��3�H;aљܟ}�N@Z�b�Q�e]+�6:�D�D,�;��2E�3 s�9^����k��k�J���	e2�����FD�׊"%1��ъ�=�O�G^0d3������	��x��Hog&�/�f�����d���U�[�	(
q�ҿnU(~�B�^I���i���W�A7G��	jd����P�ݪ%�b��b�4�P�Gx(ѵ��fnw#+�G�~Gή!}��Ա�듕��I��C� �z�3�)@�Ob�����X��0f�N�j��%��`R�j��'�&=<vVFQ^N����I������4��p�qg$倛D$(�/:��ΐ��7k ����l�����v�����o^?CW��WP޴�N�QwP�t�(�؋�Gvh(�~��&r��n$r��M��}����> �>��ɞ�������4Ͷ��T� wv뷣v�2c���#����p�E�02Q.>���� ���
g�K�Y1��-P*���z�'�x�u�H=[�����_���7��&x)�&� ��8"�bE6Y�-�h1��v:��
�A����(wD|Ml�F=����NI��Y
� l$fh,�
�ND�����qV_��E�G�&��~��l�u����
��Q4n:��a�#��E�r�b���l.��32���P�B�8X�,�5�z����n�jF��c>n�=}Z1R[E��x?��ED����`�$-��x�R���)�~Ϫ�d��E�k� x��s�0ܨC�IC#.Fpo���l.	�4�����K��t�b�I_4w�>���ą��2�I,�ہs����@�3��rJ:(�<��A�[� �����Z�D
CV�wҽn�����0+�ߐ���֓r�-~��`�~N�L�|8�o��աg|o��58��"��y�`%.�uuC�Q�>�˚���]4���F�u]2��2�f�Fɻ���t�zX_�6N�jc|�=�$���B�0m� Sؾz0���	��Y�j�QW���ځ{�l�͓�,.p�"@�L̗X��l�d�!�P�'-4w�ckha+�)>:!mQe��W��7T:a̐��a#�0��$�p��-��Ӡ.��F���k��/�}_��X2��c�q�[����z�2��O�MJ�%���2�7V!'��=�B�,Q���0h�U��z�T�����=�h�w�)" %S;�'\8��6�_Ej8p'ǌ��?���bU���aߏ�����2E����?6�3����E��RN3�,1_�#�iKfR�	$��Aت5�v����X�Cd4#�3u�k8�Gg�$f�1gO��5���8{�_�_��p�̐�NZgq\����~̮j����jH�l�T`�P5��򡜬�+��-d~�׭��@��1�Ʈ(:r�P�9�¢w���B���gG뱾����x�?%AGcJ��bc-�@*)U�����5��Z�W���{���f�t��o����cB�B&���~&�=�"�S��Q���ү�d���bX��F����m�i�,��}�<3�29>&��qc{���2�pc�5�m�̢�P�l{��k��z�*�+er�wg�~g�;ϋ����w��㦤�7�F'f���f$Xǿt�6]��h��&��R%ohU?�a���}&�8h=^�� 8���F�:�J�U�6	�8�;Y�z�Kk�������븞��uM�C�{'k3N��'���
כ:�SW���a�Ýy�+���B@�Vl�_	��dr4��C�.��e�+�n����"�|!��8 z��\:r��9a�tX��(��z��źC'bꗤ*�6T���7�XQ2}w�?�V�`�-�
o8I(����_�Qc1�Ʋ&�i�Z5X_�[?��p�L�r�R5���a�����r'�eё���-���ͷB�[��3�`���]�����H�1�ae~*!��"S�9*UW�Ͻ��-��X_���"P�mȘJ��QE������Ml�!�5���#��یR�p1��d���^�l!?PQ�]�h�yj�[%Ae��i/�^݀�3o���==�3�>��6]�o(�k������^��d�OL�^�nL��j�d�<�@��2(��g�	�F�5�̴%�8S3	H�q�L���4��?�^��� q��A���9���H���oh
�ϧFrd"WrR��(�[���
&��_�ߟ�VhX<5��ſ���"���BB���|	%M܉G���V~�d�i{J�3zo,{eZ�C;�8�](�N
��F"��;dĎe
lUi*���qQ(2"�~f^��yy0;]��$�gH�͍���(�fǔ�K��|҂�lR��v �C�����<p9l<���n�os)2e�NEȌ���*�$ڪ���)�����͆���`a-P>Z�:��#6+ld�\8�{׾�-"�8��_0G���3h�l�sY��/�|i�;A\QD���dv���)�u�P�m^�v,�ZK�������,Q��M��u��1��~g;up�o,�9���׻.a���}�j+8�����q�"���`ἓG0���Y���m�L��C�N�հ%��{�����'V�iD��C¿eU
'��/�u����Z�B9�MA�lVkh���#��i���'k�XO��J���������<oZ��4@�rSkJ�(ەn�BA�=7��B#O�n��/8vV���pӕj`�Ho�<�,����t��Z��Xn:��˚�Å�1�S?SA^�ʻ#㶎�m�~���A>��ݕ+�s2Ӓ�8ى-t��E�H��Ld�b�����l�B*=�6�`u�����?pb������_ n7�Kn_BRC�GW�@Ӯr��5�+���w��m�e���+e;�3	G����'l��D��p6{�+�6�}Py�w�����k�f���t�R�doPx30�#=���
��^����{s�(%m�����x�ި(����"T�5��k�� �-�Z��lW���r�Þ�J�z:����f��k!)�R�0�"�2=��������o��ey�����r�>���%F��lLN����侧qU�	ռq3\��dŝe���;1�'�����/��hm}���z�!B�Ȁ��+k QH�/q��G��{\m�
ز+�f����ئ��Nê�2��G����V_p�"��"��h�I����P,��gWP�cϳ�9_��@;A�*���Ҥ{�O�n��t�'x�o����������MG�}q$nxb���h��ZV�� ��
��ÇQ��r}f.���5�~JV�岆��v;-0�`*���l�-�mE�
�]h��v����a�����ٝR嗙jR�.��#�#�	�u��i0�B��]�]h��s�i͚I��]���RRU�Q�W��ز�"_���йӿ� Ά�8�':\���MY �X#�2��B�d��}�ʕ��q5آ���:A ٯv:K~Լ���)�5yʯ�y�����:Il(ܗ��L��j���ޘͿk�m��/���Ǧ/]�ZVei����^�,�E�RDwW&=�xK�8S�4D�22��9q���!mlp�Zi��z�Bf=���B'����A�K�(���c�;�B��?��sc���D����cP�d���(�{q����*��*�;B� )����;?�΂<i~46u�yj��l r30�U�A$J�ɖ�*+�?Bx��^�^�p���勉�Ǎ*�P��ˢ�}�H}+��ŕr������3o�>�"��n^���GN�K[܅��R�i� ��+�\�iO�Z!�J�<1I0D���SU�tt��\b�Bo��B� A,�C��X���}��So�B}�!���<.��r4Dm�25�J�@��ux���ua{�����OW̫��Ŗ��i��[�\�YF�t$c��gx�mv���T�"٦��w�Ȕ5FI�<}ND��.��$��Ň�dP:�&��4����Sa�SJ]i���^s�o�[��s%hR.Ns�>|ܡ��~�1��c�IE�q_�{�ƨK��W�d
W�ˀ�G��rP����D�◽�V�[q;J�R����_Az�|��%N���(Ēq��!����.�x� ,L�/H�9�ɱ���U���c������U�t�c�V�b_L}xz~�-/�R�JG��¶Z>����{�a%�`�k(�x�g�ȍ���ڒ�<�|��ZGl{�m���;�s��#��i�����=�Pv����@�#��Ca�%�8K3����E��ˊ��<T�����.Z�}���y�l�VS�tZN�p�ª��=��{�ĭ� u�o&60��]��.-�Z�sT�����9�N���ARi������N�y��Pƙ�-�����%�>\]obp�"m>���lk)��3,^��s��Ƹ>�}�ږ #�m�]����+]�Ϟ�� ÒN�iUu};�⊎y��,�OO�r]4��cBlo����u��%�e���,��(�FR���r�W�y^��fjT^�
9��0o��,�m�4`�P��:t��$P��r=i|\�j�R��j���ob6\��m��