XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���qP��Y<N#�_�˹Y��5�d-讁�y�OYl'3bt���EA80/�?2$���M�)v�ޕT����d�J���dU���_�O�$?}��i������^��rLW�W�X�u�!���IR�"o�f��gv��a}m)�[�us:W9ϙ��D5��ī$��}��'�D�|*5|���y<����\�BxuڱnF��%3ET.q�f<�j$Vy
7)4�Cs�������ԝ��Bts�|jճjd�	1pO:��-J�vW������ݰ��f����,�;�����xıƪ���Q��+ԗv�i:�DY����>�$@���̀������ɞ�>y���A�ޅ��p�'�B= ��Y"4	�MG�`Q{�������Xp<�����`o`j�����1�?2k�����j�x*�w�;���UJ����}�3>�P7�o"ζ����nqeO��c���{��f<�,��ܳ��w���۵A�j�^U�e�\ˇy�UMˎ	|ڧ��{-�~����U�Ѕ�*0�}��6��0�G�PfD���C^ya��G�����L�/W�N⸔��uzb�3� ��RS�j;<L�]7���r)0k���j0T�o�K=Fi�����G�&%UO4A�ە׸[����*C�N�q��_� ��xE�7��n�$Y5��9&��5O�
�|rN�x&.���`�qZ=:������X������Iŷ[	�N����9�7��Y?�{�J��Jjl�ח6;�����CuXlxVHYEB    fa00    26e0����_���%�ҥx���H������ �"&e�|DN.����V�o���5�z~m,tR��;:��nlu���j~|�_Wq:���gS@�� :U���ɘ�f��0�r;�C������S�,$�;���;y̯�o�&u�JJ7�,\���/��}C�S���GGE`��T�lT�MEJ�{���@�8����`V��5NP4xv#����J�0�l!�(S��B��FY+Ip���l�W��MZ�È!��y���+�����AS'��r��T�D���D�Dh{ƹ��8Ǽ�\�������7	����J�P�EM(\
��{��F�E�]�ǜ�*Q�_���D�Eև�c	��s��⦰�>A�MGu'ńxx<�T�{imA�m�9	#���=\�1�݇V���(��L�({lR(���6���+m5�q�g�sF�G*"��h��s^[-x�U@oW\ն�X���.�2S��P����`�9k��j2�n�,親�l���7=B
ƛE�ìK��{S��r���u���ͪ�.��i	�1�Xz�$��t�Dx��7���VJ��;�R��5��nd�ή�O��I0��ll�u|W����+��q�>0�O��i���Lk���@��:W`x���$]癷� �.1��hW��nꓹ?n�]$�23S����03��L�]�U$=�,�ڹ}?�a�$���]�:�%��Gp��I�4�!M�OQv �9��{����y]�8M��H$�Zĕk�̈�����r�}�-�&dզ.^ϐd �*z�����!��R�� ³���&�D�e2vw�L����x�A�����A����&�6�4F�}&Ec;����*#���c)|O= �&�O���?�cu9����5�VG�����l������?ד�o5a��5��f���]�=�N\�hPæm^���;���ǸބN����w�<=�Z��T���_����� ��D�ƍ�|^���::����q�P�y`��s#�^����w�⨤��sgiï;i=�{�N�:J�M�$�\��V��yC���W�oA�`i����Y@ �>܋�D����`��6ݛ��۠���4rW����V҉3#w-�X��MqVkVF�6���PO�K���^��'n�G���y�&!�X�uD��*8�gi%���wN��N!(�h����>1�h��~32D6��>����J�od�J�����p�"���;���tn�ε2�M��Ԯ�CQ���MEu�`�X;rX��۸��LJ�0�U�+<zq"~�1E��F�F���yf�`�ܳ�{��jX�?8x���T�in��sv
�ހ]���uK$��IcĂ,?�J�Ia�.C�8#�)��&tՇ��Fв��T0�L��
P١t�i"h���C/�t�m�|��OʌPп�y�6jZɋ���߶�~�-���>�r{�����P�:�=k�C/�:iYw�S?cfzzs�F�ѣ�Hu_|���7��wn�j�?�v�-h�٧|�ͳ��D��ɉ���*�ԣ��d��+c���V�Q2��t�	��� m��A�G1Y9��/�'��6�Л�3���T�������l�;�I�v�ǎP��1X���_흋e��bK[�ps}W�������S��|��-!���ap�6V
������o�)9.���?{�l���	�L]�f8��O���sO�Q,jn����\���h���6�ǥ�yɪi:��Z�Q����P�: ��p�R��Wk����x�Y�񿺠�`,�KM�&��5v�簨D��7$�hס����%��v��.p��>U�^����o2��X<3�-Z(C��x��7�F�u2�װ�ZZ�e��;y7�v�-�`��̸�z�e��U�R�&T��)H$�.5�Wְ�!��FUaqA�Zh���ܻ(�.�ƌ����p=���F�>@"��@�%�QϪ�<�R�4�M�4��麖t�#y��}fuF5'��z�=�%�Q$w��V�QB�����!t*Q��1������&�h>��[?9���r��َ��MR��^�)��*<g��޾DP��^�Еǒ0�ªf��B�gD� t��=�i��|(l�P�v^E�=M�ǘ��b��,��P�Z���҆�Gmھ���z|�`G:��$�Vd���\NY&���c�EH�J֯�K��ƭ0hy���tC����Y�:F%Qώ"��c'����M8`��j�-���M�Y�힣�DЛ�	]-�:�-}���He��u��XŅ4iژF9M=�v9��~J� �K�0������޼�,��-c�Y��yi0f�d���O�[�[��	�bd�_��O~�w92�Y�L�L��l7*l�.iwG�"� ւ��1���e��L�J?�Hb��H勧@�^9k���C�\�u)wS����CnWiaPZ�m�!ϔ9@֑���ҽ�W
�*$ΞG�g P�Ņ���bP�!$)X4��y����p�Շ"E�\	_1`������m�3ԡ���H�����E44��7�mcj��I�n�*��Yo�*�D5M�m���Q�^K&T�v��՛Z�(� ��!��ܗ�����G%�N�>��Fi�HM��	�r�X?Rkי}�8�Q������l�o��/Lk��X�J�N�A��)J���������j��/Q����n҉!�W��͞�L�Z#��B?2I&�����w=Z%Gf�j�j���Xc'|�
�2ѯ���>,m�'v�X{��m�/- �M�� �Ҧ�Zg��p5�_z~0
=H��MA��:��K��
� �7�>:�h�H��{�<�hO{�v�恜����c�����A\�q^G+Y��b����8U0~[8���3���Ȗ���Ί��[������;�n�.a�E�"3�V�5��rS����1 A�mw�����ʁ0.� ,����+�}KRFa��z���50�,4�����k����M�\&�Y�%rU��Է��M@����|�\c~r��3 �)���~�PB��ZR疯�'��4�N�%��T�����GӠ��Q1F0�j��qe����wB)e�������)�,7�T=w7��|��z�K_�a����_T{������*J�%�um�ns&�M����#@I�B��_/���3Ɔ�d��_���/�~Ih��1�������+J4v�~o.�����>VZ�94��r��GK�����4�3gA>�.�n�%��%f��{q���z>��L�M��ٟF����֤�y���%�/O�`Q�q�k���v��|vϑD�:&+�3��:��C?+���I�<m솱�*�2�$�+%^��T`�
�m}����"C�85u�&?�)������L0��ej��Ǿ� ����Pq�w����%	_�3���R:��f� �i7�Ϸ��8B�*=�?�ۿ�������yq��cݯ>A����o�*�	���ޓ�P�s偯fnE�9kr#�u	����f�H��VվRL���G��H����P?W�Be�ʍ�l޼����g)�}�v��߫ɫ���U
p�Gp��ΖO��P�=�yBx��@���%��Ř{'��g�������<;
��zZ+%�B��\�8pz\6��a�HQ��H�ʿ.�h܂� _*b��ESqP8$��4�Dk�d���v5�]@��������iyvk��Bu�3��U_U�����O�)����v�}��c�2�o~�������������|WjZ��y)�x�z���zv��oq����cb��$OHڕp����>/�-��=��N59�����|�$Ɉ'��R�]��7�3s/��������m��O=��2IS�О�)7��U��Љ�N����	ԅ�a\(JB6� Gp����^sbD�KT~Y>�SG�ږ��O5#X��2�9_�5���c�
E�ԇ�.�o�J��נN6�\�4��0���x�^[$��3�)���s��y��4�)x�z�;�K>̦��o��A_l��%��ޑY?[�yW$w/#�P��+��u��j=-pwZgG_o�s���ޛ_q���Ϊ@���o��(��q��Ak�%bP��f��|K_����"a;s�jly2�l�O��[�_EVM�w�_ŕMP�%_��Ax�|!aS�����{����OC��Q��t����]Ȣ��=YM���V8d2� Pe0�-�k�c?��v);�����c����z�����"vqrӉ4��mh��`�!�TU/� 7�>u���ۤv2ߊv�G+�R���� �u�n��_�]���S�^ ��F�t$eS�Ƚ����� &��3���6�CK��IIA�YZ�*Vy��H_8?:���>�T����e�Bo��� ��dvZ�"3Jb*��
��孺����v=�[}�h8�ذ�*��G;Xn��CIq��f7��]��g��Ҥ;l6j~H�Y@�	Q���t��)�p��8�f�A=�|3(*�>�oe�� �K?��hD�f;�3D;J�F1�=f�!�AEj7� v`n�k�ea�m��B��E#�6��S��l#h�sc������J3������y +t�vE0ӗ�Lp꿞��_���>�J�
�G'k�m�f��o����N`3�㳍T��ӗњX������fW�����cN^a�.����6����6��������L�f�{z+��ޞ��vT���������^�42(B���PM&��)V,	�`���r�)7��(h�}W��qM�)��2��|isY0W���4�Z-�/n�F�+�`C�=R�FR�g� 9��#&�(���� �	@�N#G�ly�e5f��I���-6a9��C��^
0������݊�#cѩV(&�[�k}���/M�a�����D��W24��O��w���:,��YcG���C�~z�k;'�i�rN2e?%M"�e��_4��(]`4gS׋G��"�1!Z��(f��\����� "a��d�]��Vo)c���5n���L�By���4�/�P�=��ZcL�ί���ͤ��;��˄Oug	j>_�@���~7���2r-�9��=0�RYZKx�3�۳�,���<J��T�ѣ* DC2�V��³�,k�ud�v�a�6�,�a�O.�#����GF���
:SQSKY*�����	��ö�s��n�hs�m��	�ꯦ�X��H7R�ޓ* ���^�yܦ��꽝[���S�yv6%���Niw�l�teC�%W��CA~�XB7P}�5�)�V���{���� ���(Җ���'�����)�4	���9��pjr�P��p��[�c �����ω`�ͤo�X���Q�w+�?УX{�����(�=�HR�:�ޚѶ�m!3����O��G���W�/���K��	@��\c�����lK�Wq��S�CDY�-�˵���z'��.6�uwD��\߼6�\cp��_d'�4&��e�
D.�rF��㔹�zU�Fn >L~���2�ً��DT^6.���r�ja9�գ�_����Œe.V��ő���c��m�B6Μ.�ئK�>{�<X!���ʺb�O�(���2���	����`�F�37(?|�z��a��HJ�0t��^�ב2x���'샿���"�������f�c�1\ Mx`���|�=�3�woU���}b�3�b�������V��Ou+6�<��/�ʳf0�d�`ydR������ O�*u�o��4�O��HU[>mB��zh�ٳVg6[��KX��]���Ƕ\bfŅ^�1z#��G�E�}��p���gb�Q�ht�:P��-G��m����.x����r�ӉdMC_��)�f�t�W^b�eS��T���!��3j������X1N5/�@A1lN��O��� �;�5Ȑ��7	�W>ɝI�%���(yu�&�[��M~7 {�oՆn̹j���$�z�����	�o�6�IzF���w1�Ӎgòt��qò���d%�JE�4��8`��۪E�m��'���RAyH�y�k�6�O�)��#TG��a��-��ONd��]��@�9f��x�#�W�ǟx��;EW�B7��|�V�+BOD[�3d�Y�l���>�)8K� ܅D�vu"��$8�QN�fT�c�c�$�U1�I���œ��;���w��^0���/����&��t��iTu��,�X]܈���^�KK�u9y����iٱ?T!�Q�(	�I��U�į\ш�Đq'�q�)o/Y�Y�}96�>[��K�'1r��Ig��}��0���h�j��K��<�#eR��;���z�^˟�^w�����@�����B�+Q�Uj�P�O�X�(~���3]� @n�-_7Zp���6#Sty�^=#I߾��������g��(�X�-�����oN������=�'�uq��,mHX�p�Gw����G�~5r��ܮ;*IGXK��������DA м��$��P)������N��2�طmp��k�JO�G��9���~�|�����7̎}�k���m;C�PL��ɓ`T�]��v@rD�;�Ss���*���d�
�]�	lM=K���S�-���ߞ�����#�3�h�ƯVA�ǟI��"}\R�-���.^��=PA�_����h��ksu�����63��>�9�Wq�JQ:��q��dιp� �62��i4���#P�'��.!��v�{j3���sgթ��K�/�H�s����:�*�{|��}������-���)_O̘�,#M��y1إ���<��!��{�Z�ʹl�?�F�i5�5�FRa
��O�P�����lN
R�√AƝ�s}2��@��=(sx�rZ�J����U�c\�\R7���`' �*�i�]s]����r9�7f��8���#�������vP�%��#-�ZN��G��W���J)��(	�.�e�(�ݏ�&6���=f��T�&�fۆ�C#q<0��R��2Q��* �&��\�'IJ�lC���1nک��v:O�^�c�qҒR�5IN`��l��2�g�((��V�-6qh��:�AD{�Y��C��ͣq���h��o�����sp�qύt�e)T����t⼮`�_��f�~K���|L��'g����j��fy�8���\Xk5  ���f!Gde')��~��Ey0`"�~�3�J�s�'����BYO�h�,���(�mэcҿ�c�q�x�&��UU:�˯��pߟqFp�*��o�*�2=Z[ g���+ۋ|ƒrL���=n�#�9.&-6d���ZW�D������giҎ��k7b���=+8m��p�"�d��+����uh޷��+��5��\;����xt	���"�/!?�EQ�0}��F�4�K��O:\�ůթ�$\�(��?����j�Hf�߇�x�šr��� �w���"��I��閍���ݎ�0�Q���}(y��m"-��s�Y�vN+.<�:ۜ)jX;m���N��m0 ����/id�A�g���5؟�av���E�b1�"����T�eX-L���ځs& �ވLj&��^��A݊kr���s����E�;�Y��r�C�Y���A����ح��8�ֶ<'-�0�&��	;���?%]<�_	���L6ؠg6*Ŵ`��wCO<H�M�W�`?�%r�X�8-i�+�]�&F�dR|���bU���d@�YM�H��@��ӡ���Ϊ��ps�.$�pAH��(nV�t�m��j���]�PM����#o�[9q�/A�2Ps���F���G~���#�Y�Q�
}
��`r�m'������S�W�eT�lG�� T�)�D����n�Þi�����ހ�}��y��a�afEX��q�+�c$ذ<�q)EP��`�|�E��f�9�a �Qq��#vo5l�Ie�E&����=:s3#k�Z���'���bS�w2TҚh��@�"��rL���2v���>$1"�]7�b������**�w�͸��� T'�����<{�q8�h�Y��7%ߌ�C��gC��Wn��>K�5���|*�d'�����J]f!t�띌�<�RJ���*�� 3����M�n?��|
���0�2 -�?2����	�Cb���9�[���~�:���y���:ͤ�Ǯӗ�f��:���W�;�'/Q�%�7�C��R䣥)
W��Y8s�N����r	�/u5HϪ'�#O=�Iu�d��#��!�S��&�w��/�|
B@(��)�l��]����bh1���b/H���iG�-R�$	v�BX�^����j����y*��|�l����~h%���edcyV!��Ƀ��Ҁy��܏��T�)�OUPR6S��Y�@�g����g��sمrM=��kwx	�n��4��	�+w�l�h ��d�A�x�N���/�E2a��ܳ�}�e?���F���S�5Q��_($�iզ"��h.��y��Ȼ�R�|��O��D�%�Ds��_g>��8�d�A�^���[�v}�T�;�@�`��W@�2��E[�5n �hO����x���X����y��!a_��_�g5ke��'����I��؛�b�=b��pŌ���1Ahx���0hK�?�XQ�.-��J�gA���3�'�.�*{|12Sٶ�n��zb$W����{VTNf�4�=�Z�����Y� �<���GQ��T�{\�_��g�B�����_~}�n�������3pY@NGQ����
/�T
r#�#Y����M�?#uw�����Td'��N��݁Dy���|��I���0J�n�����A�����H�s��d
<�Tz��+i��D�>veJ��B.�!�J� �P6:�ʝ*w��	�@�Bl����b�u������x�o>�N���r��)I(Mj�P��'v@&�{O�ھGX��x�>�c���	N鲀��K��Ɍ���Q::y�>�chs��io�{QĞ�Ρh�4X���'�Gqݿ���aem���e�ړL�e'}����w5�"��?��9�JN��̎Ge.T�)˖�����d���a���Ry��$�MP��7���=i\�me6�L��/�Ķ���lȖJ��pL��/ͻ�ɇ��2���ٸ�������&h��zS�������j#��Y�}� ���]��w��D�G�E���x���V�n�P����H+���C{��z�)�R�åɐ�*���β�Y�l��S���v5��� u�=Ybj�h1�1�׬�ם���T׍$�52o�0�V�w��-&GA�1��	N���<�������|�^�}����C6x@��G��R�6�47b��O7P�$�n)�I�o2�qi�~(LD����ɵj��=��*gtk���m!�:�m��すJM���l����Tx�:;�#T`���+jZ��q3�Q�/��֨��>,R���]�Z�yk�v��;5��+B�%�0��PD����D{E����ˉ|Xe����BA�V88_@vs�b��.6��K�We���U�4~��J���{�G�uIN뷮MI�4N��P��"l�0�n�o��(�3]Q��)b�~�c?�QG��$���Kc�G�'��ԾVQ�8����Rش�◿)(�����p�*��С�$����KN4n�����O���N�rί�UJ��]).כ��\g���b��>^8tۮV��F8ŝ�׃u� S�Y��l��6����z�;-N�;�3����MM��T�׀4��^�ouNI"�I���V�-�w��3j�p4�y�"��&;(Gٝu�¼,�Z꺚���`;
d`����X��}�d���g����ӄjC�jp��3�ㅾ/���leÙ��/���C���,�7�)v��XlxVHYEB    7d55    1450��e��^���@gj&sVc[�.�g��c�5혫=r��Dib`s�8dJ>/��b��/������7�:~�)9h=�fԁ�!�M�/��dQ��Aab�(����V����d��<MbB�6-g�We'�WF{��[�_�U!���4��=��j������u�it11v�ҷ��;Y ����e؉m��P�h�w�$*�LDi|�z�ϻH۹ѝV��	f1�O���"��r�o?#N�#�m���w.<!Kı�U{H���A�q1�(Y~�j�}�.2��3�Ҹ���a�(��3�gEh-�¿�r�fo��"��00t��6�����\�^�X�*�^�����%]P������N��I��_�6�'����/_����F_�s�w�Xj�ҋ�7಑lu!l��Sm�Y϶k;ʧB��ҕ��gx�h�D�m$ږ5�N�V�����d�[DcI��f���=b\H�㍵z��8ٰ
6��m:$_S�_�JC�=���\�C$%/��@7�u�	�����m�FP��)���ǲ��Z/��L�' �0SR�Q����%��g�1.߻��m�
U�G�Xz;�*
W��z��B�{�̮Q��a���`\O�NR8��9R5\�n����A>������g�)��H?=�V�l�'�ˇkTb�o�.@!_�g�S!�RU��job?t��Q�����+G~ �a�AE_o�?<@I�2��Fۋ�j�v�H*�p�.�x�̓
a @݁"�=DNY�n!�Ti�o�Ҵ���]��"�Ua��x�U48!��\�;�]�}B�Q��Z�E����:�P>Sf!���Pm0f6�)�&�5m1�y���Ѹ@=���N�Le���~�e�W� rҸz����-�.�^�nŞ�a�ۚ�jG1 v�ֹ(gJMZ�)� ��ҝ-�D���@P����YZ�o-Q�igQ9�	� ��;��L��4&YsJ�B@cl�=�,>���
��4�g�F�
%,��- �`��U��j���)��f�z�~͉;#*.�]��>�ؓ�V�֯����Xw'I+�����|K�(�j9�j0��U�������P#�Ζ���!��	��v��	��������`m�ԯ7�v5����!�U�����t@`�ؐ̏��2~݉($��4��l!�������� �sN���j�:"��&1�ѽ�A���ĲӊO�Zn��G�U/e���L>��f۰�� 
��A'|b���U�W���;��	�i���p&J'��@��{��8T}g���27�}@6��H���26��57F*��5��¼׊��a�Hh�o����W�J�U�-���HߌN�F⽸֝u%�,p���,BA-xxuaǊ��n~��{C�}�	HyV����Cy�á5��R+鴅�̴9�t�ƚ�+Ȗ�����G���$=�o7�G�����8ԏ��nM���LVL�þ͋)X�F~��p���~3u��I�t �����x���h0��0��j1���Y�����O.�1Í./�Ή6�5�S�d!�����t$�s�3$1@.S,�F�~�u��@��2{0J�8��*�x�6ѿdh�����'�3⤦�e��dF�����-�+/�2\ln�$�w�HH�����Ue�/�]-<���!C<U��l:��U"t�f3� K����ݙ��U�8�p3R3�d`#���-�m�q�6����bl��&��Q��Rh�C6B�%ʣ��`���ŀ������MN-sW�+!́�������i<w���UY,�)^�n��3n�A��8��<LS�LXiw2���D�� ����}G�����w�[2��e��,�������m;���y*��߹��
�:U2����h9� �#����YT��zf2�</�3U�x�:'e��|#=���������r�qK�8�d;pL����}`Z�C@z�XB����s����7C��8�X�g2�{���~|�ͣa�{^�K�a��q��4L8��
�b$�ж(�&�l��S�m?�����},�n�B�����X{L�'x�MBH�Uc�펴ޜ������`	�f��L1����/N8�=R�y{
|=A�Z�{!; f����e��6>���
�];a��ۮ�]NNf/����
+���`���z�$'�0| _}���aat�E��`Ԧ�Y����L�"���Ko���џ�����~��v��{AE�������}+�kZ�$gZ��b��� %�����g�{0� ��/8膽`�¶�@��dԽV����T1�5��v�!�MjGd��:���^P R�����(��I�z�`��"�]�h�*�}v�>_z ���Oz��\�\.[�a�r�����*��<�N�?N9���j�3͞4��m������8�j��s�
U�:#����C��zP�M.+/f�4�Tދx���N�Gf��p]��m�AɄ�*��rӨ�M="4��A��  &�v�����_o�<�����
���[��NՎ�Q?�:[���a���	_��W(]،��,� �Em��ǚYP��S�޵m<Yy��g"S���o�j��Kؓ}�a�O����]7gV��.z�CA�����04��H[|[*�}+JA��?���d�:��5	�m���z����%V%XCx?S���\��?6PFx?�&��F}��H�{��Аmvv�f7���A�号߀�[��c�Y-� �:?Q�*��3�r�f�{�<���L�O���;>3ܞ��.�E R�����|xSzYIR�K�զ�8H�u���w���A��;�Ȗd�l�M6�2�of�� G�:=h��e�v�;1�9e�����oV��.�Z7D	*�W4���|ϣ�
)���_�l��Y1#X�h��/0���N3),$�T����tq����lfD`��7Q�Oq�K���r�4>ŨEij�~��l�`�#�;�FM���t��?�c���~������2��u���wȟe0���M�)N��ԗa�B��lZi�_��Suݙ���-����]��-�F�鮞c� ���'�V�4���ނ��Z�� @���q7C%#ig�� L�2��ms���М�m��9�?��08��Z�L�MTJ@h8�#��0����U]��g�U=�	E��wH[ya�_?a!N��K��<���R�z7W�E�JU�����3�?ֳ#�yB�(~�=��F����X�;Q��(�G�5�ƚv�J���wō�8tO��ӛu�nZ�a&'�{��p9��'V��?u١����gn��� ���z�:f��8���*���s��
���AX<���kإ��Y�4؛�¢	�I�@�s �����cm�ͤ.ne�>-ˤ]ٝ.
P�c��5>�21e5<+�-M�L1�`��v
�Y�	�h$������LW�\>V������OS�^�e�F[���a9��8���N�������\�$� ���� ����\���H9V1�v-%C��'�f�ao�ĸ��3�^5��g�,By(iX�q��D?� ����B����V�.�"���r�.��0��'w��8#u&�?ӱ����e�:��C�,���?�ɜi���/l��;M�8%�x�%)ȵ}i(h ����R��c&��#�UK���1-v��4�Z���O^�H�Cf�ܪ6��	�LwHZ�܄}d\��w�Kp��cC��IT�(1���]�3��zb�U�h�ER��Y�������'->U?{
��)�Aaj�|I������g1,��#C���G���x��g�	�R���stW���Lb��9�{O�Y��Ny��=���%+��E{o����m[��<U_�5���S��j��['x]W�[�����#�iI���y�Qnf�!(���gin�(�s�\"r�P��4���x�B\�uM�8�<�KO#[�.ꛉ�B-�"����5p��O�ܪ[�r%� ��|9PѤ��1Q���L�H�����1��Ha��h�LPҎkLͨ�̰�2�)"rҐ���,��c1�Hj~�
�ѝ�-j�"$bp�� N�����j2��=�����M���캑T�����5clw���K�̪��4b�o���8� ��%��hv���a�j���,|)�Pl��Q*��p㯜�3ҡ�_|0{J`�?��foǩ�[�[��>��G��S�⏂!Gf��+�,!�Dٙ�$�ѨMR�;����q�f�9�clZ�N��l��04o�Y`CLI�sm�lGb��dV�&�}+
���a̎к]�	&��{�OF:�� @�JY:s��9?MT�5�(���o,jv�r�W�� oƔJ2e�$�_<�q���'H�şCP���ޠ�_�_.���9�f;�d�.%��(�T�y�}����N���)7߃�����B ��'��G�<ɪo�ۉ�%^�E5Vf��_�8|*N��U�,�ʙ\6�+r�I��O��v�
�sP1��K�' u�;P�p��(�'IJp�u���5nh����LjkOH�BЈb6~.�q0,�H�����u/Wч��eu_�9 �R�M��N����B�4ð4��>#l��X�lݡ��.C�V�ғ�3]�o��g�"�v�I5g�0>&6�_�U]D�Kþ�m!��q���Uj�Z�;9���G��_m����Cn���Ǆ^e� C3�Hv�v��ْ�BtNT�P)�L��=���� �YM��2@��E�k�A!v����9��z�ӏ>+�@�T�暯Ԑ�r�P�����$E��V��d!%�|+ EX�I�v���)�o��ݒ<����ָ-���i�iūLb�}1�'����\�]KXݸ}+b#�������6��!M�*n������;}�]��j��d�f��xK�>���IiD�ZL�D�����T��<7�|�N��;kX�0\џ�|��b�Z��|���>(4�jcs�`h�p���pd�W��h�
��~�-)����6Ө���M?HyX-���D�&g͎
b�U4s�c"6�ɴ�8`�rcu.<����>�^�Z4�3�͋��T+6�{�j��X���UNpO�x=V�/�dpf�,�;X��憽wL��_�F+��  �T����g6,��w��e��H̪/��9���y�^E�'!�琓�ﰓ��|��7�F"@S�n�~�