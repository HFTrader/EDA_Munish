XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4?I%�%�h����NpU�2���d�sg��~��A�z:�b�%Z5v�Υb�>��F8�ݮ�m���K�S̊؃]��&f|����8����u
?�~iQm�޵��7����<ەJL߿(Zc�b�=�	���E̓ �l�K[ޅ��&$st�Ve��3���e�q���uܡ�:R�nOe��^p,y���V_I�@}y�ȶt�?PUf���
��s*Mfw�J�"�-��ɸ0�rz��U$�>��8aCy��L���x,���l����~�����<�0���2�)o^ Q6�di�5G� �z�E�x)���ucf�ln~$�t�W������^ �<l�Nii�QL}�j<��o.��F-|J���P'b����&��4�Ӂ<:8P�Ѐa����m��??>���Rp��`*ď;t@�=!Y��</���9�P@|�����L<��(%�[6������^��1&̘M�
����-݀��"��7A��3��^DEis��1)����*Y����X��!�hj�s�^ʹ	����j�|h=R�ݦg�Q�|e�aQ-��˨�]��%B���Ȩ~����t��7^-��i(Z�=.`�@<ms7�ǎ������ζ q�Nl6�7�P������p�&�M�ȳ��<{[�R�0�-g+E��+� � I@�Y�@��[H�"��{�O��F����4m�M@X �A2�lm]��/WLa���;� ���ĩ����!d�G����p�-q���(i�_��V��XlxVHYEB    fa00    2910���1!��xx"G`}oA�S���a,V�$��{���ჀBH0�*	k�LV!�w;���ۊ�i7r����F�M�a�ɟ�"�a� #7�q���H�&�wZG��&���+*=a�=�D��ԫa�v<l�ay�R<��M�J�x�&�ҽ8GR�}s��>���H�
TW-��TH�x�T�*�/:L�*��ei��S�a�(�G������/]W6e��4���D9K$�	�p��>mN3�����A`��Y#m=)'��+��f᝻�$��;������D��S
pV�*J���r��L����N]p�
�Q/i*s�β܍�U�wC	��1�Jߊ^պ^�,E�����AtBK]|ÊT���i����d%�l�:��	���OT������:	��L27�ڀ�&�ZM��2��N����jꛭ:���������G.�n�R��M�wRw�X>_��q�y�y�`�Ub�7Y�K���V�1��5\�59���4��Y�.l9�x��IIi�	fr��a����j�~ZB�X�ל�0�T����W��&}�_�*7' ����Do��[�o�TU���}���jc#ɟ"	֧�IPi�A�o�u�m�/7h%.s��SlL��7��CvY�j,��!�p5~sQ�8�͛_�^{Us)��a�.�U�kuqde�R�g�����l��~�6uƖ����>�B�W���IS�J�>0����c��$IIj]���y�tS���9K?�u���`���ʜV6����fܑ�rHT�X���cex+VB%��N�v�6۷�
\�M������ք�4{�@p
�K�r��K-�(����P1�?�)�ш���]��R���Đ88H�a˄k�a�6�Z��I���i/�\��Ե7{T�����F� ��+����s�==g���;]�LTW����R����?v(�`��_iaW�|~wk�4�"Ι�x6=�ﰶE��I���.7\x.]7�Ev�
f�b����u�aco��;�j5��ܖP��K'�2�p���OEN3!Γ����OO�+�rL��;ۀ��@�(ؐؕM锜s`�Cla�Cr�:�-��Yǝ���f}��V0 ��5;�c�����Cn�噀&�vA��@����<gQ���b���u�	B�A�s�2k���Їcb4E���N�+or���1*���c�!�_J��B{e�hN��l.��?I�w�Z⫧WǕ������H�.]pE��$V�}�)7�����<��>��A�ٗ�L�Rcw��3�fQZ��i�=�b�F�V�?�HZ�0�
t�����̤�|G J�GN�ߪ���9���
��q�W�����M--�[^����]��-��ߖ�
�2���_~������� �%ى6Kј��B�� ���l!��`J�=Z���V��J�����e�����?N~d=M�c �E��Ms)?��5Y�]��U����\��� Yi��eO� ��$�.�HC���R�+�H
��E^M��@�f>�1�g�&�6t����"<4 �N���ӱ�A�WrQc�j�}5O_s��{�:k_��I�kӀ��4H}���e$�vM&@{�����!t�0o�;�d!����|(0���n�N��>.�ͧ��x{b����7(<Xj��m�'�F��M��Kt����p��"U!,�:n-�PdY{2� ��8��{����;>.�9�����3Uoj2�7�t��,�pE���TA��<2\t�\W}i��m���C`���*�hG��$� TFR#��/Өå��[�b]�ћ�q�����؊���c��$k� �n�|���[�R�[�/*�KV���h�h7X�9v�$�ʠz�a�����x;��Ux���4��߫"��oGY:�*4rV2�������ʹn��	e�����OJ&�N������u��4���n�'d��_��M��9�VfY)�k4݉���|�E���"$�i�����0��i�tc�bZ��|kf��͏A.Q	��-88�D�D��3�)�OWC����'W�'R}^߄�ĩ�������th-?�+���	Iy��oy�2��&3�X�z�)7`\V{��5����\3��Z�>�}D@h���I�񖌳�U`n�"���@>���:S�u�-�E͑.a^�\�0�8��vh���J\��?�A�@�|I*�{�����/�^ XX7��̀�8eak�7��ErB��f8t���j��A�-�z�����CX����*jF,h4σ��4r2!��2+zAn@?n�	�.��n�q5��ܲM�� ��@�t܌" ��b�>����,�P�̦���nw�SWV��~��ņ0�)��X�V��6$-��/R�&i�W�$�K\�/ ���Nw #�;ɆF��5�n�v��!S��J�,� �,��D��C��ڄ||:7�k� ɷ�L�F�;�2_\��[�j[I6��WS����T���k=jӲ�����j��4r�׮�5�p:&]i[��"K6(}_�ʇHe��j\�"�-�}�r���0P�&�����g[!(~۵�+xd�m��̒Q�T��B�B��o�C���ʖ���܏��,iȕ��O�Gw9^����V�	x��!���L�:�n6�[���i�ƥ~�`&q��B<Az��&�T����e���	o��L�GN@	��o��X�п��
����W���|�$.l/"ޒ����ڸ$#F`��^�������־)�ι�΢���rc�9�C�?C���O���Ś�!ӫ_d<1mC{6�D�F[��"��^�7{��R�Ì��ZIb�ɼ� "Zv3��nF5�:k�t����T8�W
��d2 x�L�2x�/>%�f���@�&�o�`�.�?��/CB�:��5��ah5����[��>��CJ�Ӳa���L`=Mȳ����Q#�; 6�q��3+��p�׶A��w���6K1;�7S7�ع���F:� ����IX^��'�ʧ�A��*��𓽇J%�}�"�u�:�o��DC�w/�^}<�(Z��ꉪG,��x�4ԋt��Y>K�&�õ`�Ƕ���LXZ��t$�1��\�-}�$�8f���g��P�)���(<"!��?��X��~<�a������S!�����!3�tK6���ۧJ�VC��62�jh;��:�} �@�?mA�H@R��"cм1��i�Rt@�%z��XH' ��n�K��	�Y>t�#��)�� �K-���a�|�p1�a?u�o)j˅���.��@�{3�I�#Ev5U(�=҄m��ltyVKr֝�Uq��FJ�� Ҿ����{�k>�PPr�J�nm�Ve\��Ӊ\��/�"-�oL�Ug�w��Ьw�SY�X��>�W�Z�9�H��Wq��`R\�Sl�a JhgX8(���.�>�]H}5�=�<�n�Ǐ�@H��W��G]_a�$�����rsǯ���}�5���Y���_t���W	��L1�̎'g��A�D�2uy�����ؖ��w|�}��I금�w	���P�p��<�*)|�=E�>1��͚w{��2��w.h6���o	��o��4��V�	U/��|�Bn�#h̿z�/�M�IUq�^k��c��,��J6����X�y߄:a�ߦk�V/1cW��@�jıdN���=~}���tW�}�����H'������		�c��'�#�b�rZ,��u�U+���No�M)���&x{�= ��M�lx�MN�y�II���C ��-I��{��]6{��C�rZμ�x7	�h���� �O>� ![R�9P��
�6���u�=M���w$(��B���+���xqh���.n��Y/]F�p��'_��{��\R��(�7�$���(LF� Ε�eFin=2^���]*�i���	׺�uѧC��P�ͬ/IgU&�ɍ��n��qa�#�x��;�s�i�Z"/�I��B�k2���0v���@@<BrE-<5�d6�E��P��`�W�}=7����9V��EER�<f����+�2��C>�&�<*�M��<�$��S�+�{8bD����F�e:��kE��u'D2�μZ�twŴ5�&�Ң҄�v]�|r�����+՚n�~)k����b�7�s#\�����k��:�%�!Dst
��Kz�ߢR�����p�����#���ЦV�ʸS����8�K�jkڤ)��}-�^Hb�������O��"Kn���rqs%�������Q��Kt+�&���\�!�d;B#�3�0��~z���&-YgR��$DSxE�*�������s�x����􃳵����X&��
�ف��gcK�/i]h6k83L`F��؏@Z� �]���V��Г&`d[?a�M��mZg�*k�	�Oz5lbo����aρx�U�T^;ED-���X�9n[�q���?���o��;[�V����E�ƌ�x�J֢6'�z���
|�laP&�X?m1P��/��8��}����e���Z5�e� ��Lg�7A'bz��NJ����Y�-aT��J����<:�X�*+��������څ_G�#���6���TJʾ��ҕ�	�}�u��2���U+t/8�W-�A}���@Ñ1:N^�K*.L����f#X�E���m�;1ªt��=[F+�u�>�L���̑�x}��bS3�Ŏ�	㢳ʢ�
ז�~f憭�S���C�=;�D��� rDO���-4(+���b��iy�2�o��N��#��5I�.�&��� �$�.H���R��|���z�C쥐m��~� �	P��	�*�R�� SƜY�]��������h<UvB�Gl=Xʙ��C��-Jd�8r��1�.��n�|K��HQ$q�=@fH�**�>��+��f�%�k���b�i�6YS�+T����Ο�S/� �Xa�E��J�pH#ԄF��eՅ�DaSl3��[�Tm����G%�y].'y�YdO��!��'�����rR���W��/����2"{���:�}�7���{��u4�%��)4*��c@���� ����T����q%r�ꫛm�@�ekEYr���̻:{2�Ye��
�!wW�]�f'�#]�Ԩ�,��!LGQ)�]^q�w����
5��F烾�~�t����F{�g�z������;����4)c������?�"��Z�:o���
��$�O
kq�OΎ�ݡ3y�Jr!j.�xn�zm6�=4C��`T���t7�YH'L��h�W��/.��4nc"�������MV%�X4��kf£�:��Y���fr'u�/��a��w(0E~�n��>��=���I:H��(�@�Z�T��ߩ6��QI:1���%'�~���K�&��]!b��>D�ρ3���~=l�`>��w���q�p��eDydB�Z����?�~h��)۞�ؕ0���~j��5�U��z�D��<Y��k�g�}� <[_��ד��Q�	tk���ٸ+Q�U)@�H�7C�uȹ� mJH�'�ìM�q8^r���ې��?~�kˆ�*��Ea�~�Q&�����~|�X��s��ר�c`��Ċ�<�//�D�^���6/7�_��5��H�&+��w�CF�O�hS ��:][|#�|����iջ���"m��]���3l�d�~߀L*�J �Ė��E]�o|`�o����F���;G�M�s�����4p6�Y�+N��d-�����1�.�?X+�H ��ኲ'�Ζ�J=U�TB��
ʖ�(LG�N�:��_Y���bd�%�޼���/_�S�����'�2��^�@�4�,����U�������1m��w�g���^ۛs:��
0��Jǵ�W K��y�f,�E���̿�C�zZc��+\���|x8��?C{c18�}�Z�#��o�ß�lg.�Z~C�;��s n��l�u,����C��?c(��ف]2,m�.�/k|��蠽"(�'Գ�]�����8A�(�����i+}[�˜����*۠��R��3�O�d��%��][�B��ۡ��2�%s��P�wy���֪r�"�d�/� ��_&�!(�+��;�A�Y1�^���@�{�S��R,{kdZ��a`�����h,��(qW�n���s��V+�s.�B�P�K��hsNH'�\qf��,,`"h��A��![7�ɿ��+˳)��2��0��.�H�j]��i�	�l���l�Ly6z9�/[��T��eQИBds@+��$j^z�ފ��vfX�@[k���gѡ�?���D�u�X<3��_!���[m��}mS�ގ�}D���d�\K���H���B��;����ۯlg�_��Rv��Ê����G��@��v�I�߶-.
�:眪Tc.C���!�a��!\��%|�JY�Z��LpԴ����0b�P��a�>�=G�M?)j�IZ��p 9G���Rh��xV$� &�0�����60�˰����Zf�"�3�tCRd��>/�d�0�閯���]E��p{�Q
��$�A�8m	�=u��S�}�^�2r�28a�P8�&�n�g���oi�^! �j���`v1�L��K��	0�����ʔ�a �$>Vp�͟��l���� �Z�A�H>�74��b�a0"[�����j���c�	�=p�/s�� 5��C6��Zf�v�b�&eS	�y1����X���(�9њ%�|y���wp��/4�K��J�l�#������i�~ ��?Bb��U��Lv-�N����gF�'�j�{�Y�������D_Lyֲ�Pd���g�φ��*�{�?e�\�
N����P�í?��#�cw���T� ���������O��~HS��r�#�B*�a*��h:v�n����y�T>8��sU��0<N@�f"�̯�XY0X�/Q��GJN(��FKª�W�	h�=��tʵ�Z�����jו��ꑯ�O<��^���ߍ��U"e��4�y�5��N��"<N|�<e�\��̭��	�Ct�����
Yc>>1�MLax�/���'���J����,;����O��(��Dy{�,C@�5�>(Ҡ��}�m����KO���$�;���2��NWԠR�;y�FȬӧ�*S+��E��UZ�"Ƨ7��Ho$�Gi��S�dϙ�E����=²`�k� ø�8R�(^_P��ܕ���4�A����^�X2*�nYY�g~4X� ��!v���<qDWc������%#o����D6�%�ņ�&�r��0�I%���^U:$��;�H�y���2\�[�͝�ƸQ�>�R�r��b$�e.��$���Y��4Y���y%��+u�$)�X6���6���������k��������o݈n�FI^�1�;֨>�.�=�m�M:(��7��-����:����N ��6f�7r�~Df��1���L!��*\ƶ�A�Z?�A�1C�`S��6�"�X��1��_ʋʣ�;�}C�b	���5A�T(Ȩ����.7�MM�C��l����_1@\]R�)
��n��*��B��&-��j��s�K'��<2W�E�	XJ�펔��j���W�sD�=��J��o^P�:�,_��s�ض=�:�A><�'d�z�� [g��겇�߹ú�W�<�n����côt���G�$B|^v��w�0?ɚ��*��Й.��CC�J�.���y|l��C/��h�21��B�x���-�F�*�Lw
�J�>��W��,�v�xܮxg�4 �� յ��1.D�(�~��$5�ҹ�bz��5�MJN�e���7_��$gSs��*w�?$�����&�Ҁ�2�C�D�����~3�Ou��]Tg���ţ T��RRjqC���f�[HMpyC���2*�vEū��萊H��J��Y뽛�w(�����]�d����8Lc3�]}g&����r	̣�a��q�8�k\ƈ�8��t'x�@d���$(n]�PovfmB�88O<�uLc�h�K��]@\��#P�zއ���¤h﷏���f����]͆������l�o�SQߦk,��w՝�^�X=��H�C�^
�ލu��e�d��a�
���͠�		�]�y�"����y6L8�:c�DU2n�Z�L�^�2R'MK�)���u��[_>����em��S�J��^z�7d��#=UA�>�w�z�����3�V��n�65��#ɦ�!��q:�!T
��:Xq?W���mu������ ])h�?F�%B x���/aǴ,{N]��b@X���w���'��X���0%y��фnX��Pv���ą-	�w�@��[aҗ��n��~�wf�-,�!U^���
��ps��:�ջ�э>ZN� ���:D�<�x�e��->���r��!RA���d��y��|�!�f��;��5,����'h�.^
KVr�������aC�_`��)�b�:*; �c�pih݄7� �����a���w5�l��W�@�|x���# u�5�F^�� �����J��x�q-˚��W�f��l��O3�WOx	n��������|���G�Una��]��\I�����3K�^�ߞ~pך�+|��³�iљ]� E��b単c�\�Nd�Q��� �'L�_��?���0�w,c:̬����ǭpB~L-6u�����N�"1��J��uF��Ym��Kqӟ���%O�$�Go����_㒳�|/V�������p���$��'���m����R��[r7ϻ�)3��P�e(d���ͬ�:L�z��w�A1��KG�DKn� "-�m�V}�V�����=�h��U� �`�JsZe�_�G�I���z�S���/��p赛X�D6V}��Fٹ�)��Mu4x}��#k�H��LS
��|����@�+��¹) +�q\�b^muGt�B�U����Vg�j���B��r�h�{�O�=|#�ݝ��'gf�U�K��1��h���(-ǧ%)��ƴ����w���{RY۩�фh����*-�[Wu�ʒ#��E��C�jdD��q�'$�P+V�ݬ�ҞZ1�6�Y@'�c�<�}�MbR��]�Z��B��%N��غ�§&#�́L��J��x8�~<���F�BHXڪ���6�yl&&�ZB�c�C���:�:f"�����H���.�/X�0������x$%c�H�ij�-�XFl?0�
�#�L�9�^�0Sgi~2H�0j�6�.q�#������f����E5o8�Y�W�����ص,h9�S�+4/N/����^���,��~�jP*�\0���	�5O΀� O� lo�����LG�5~�6��O�2�G�
T�g��\�l�@����`��|a,A��@�
ir\��l)W笪n�f��.��/�G~��rJ#��Fx��mE�j4��(�r*h��4^�?�C�.|*��V6s�EnyGg�������g�ߞ�eKWV� Y������}�LxX�qw)z5��mY�FZ�>Tl�7��ުgѤ_|
}s<���&�A�v5����}�b�f�jV�gWC�5A C��b
y�U�����/M�s_�)��O�ܲG5Y�������Rr:�w{��n���|kv�Ѻ��l>�훠V�LGak�j�	��P�Q~�,ө:9X�/�K�i�m8�m�
nك�B��S��9�F��Ď�_Q���~U�ɤx��k`�.��GЄ\% zan���D���΀}����x�F�/�f�"���������Ea�B�<�:�D�:�{��d}� 2���0'�qK���ͻx�9ַ^}�_k�=��N���P|��>�1����Q#	��7�����Rx%�c�PJ٥*���5ˈʄ����J�ٙt�Y���㑆ͭ�����ﲷ���h�{�n��J8���|�=��O���T�q��x��T񸻓ۄ{��g2�sHy�-y�`o刕џ���J��|4rI�Y�<�rء�b�L�a�����7�q�/�A�[U�!���[Q�6\Fo`�0���SFb���E�~�<0��+|���8�>o!������9`��g@aD[�	> P��>N:�aQ?e� ��.7�ڶ���b��pE��h�&�َ��.�ű ��Am�6v�B����d�/��Y=?���:I+�p(Wg�e
�Ee\mD��ð��*cW�
^x�$�IZ�7�|E�18*Z�J�+���/�&, �%�%���W����L��=�
�b9̺�$���H�u���N����ߋ >[Q�ZSn#U28�b9p)D�vR�4�D���Ŀ�N��=3=������h�D`S���Rqx�@���j�кu%s����=Z�����(��dV��e.ܜ�c���������:q��[�w϶	���ؗ��Bu}A8�5t�:ս)P��W�W�K�)zRa�Ym�	8��̙ߜ�/���q���A�Ʒ�`l�� �h6�Ө?���u�An�XlxVHYEB    fa00    1d80�phzm�����+/�S�`ޓ��a2��j�>���ʙ�3u��#U2ߓʃ"<���K��̦=�:��w��;�(���2L�ݛ\���cZe�*�gafF�FI}��ǛH�^K̥bo��I|Xy�*pb�P�$f�p7���Q�� q��;J	VM��ᓬN�b
��B�8�f�N���C��e��X	0���H8o�>"�[��I�ZL~���ӁkO;'�Ҋ�"�;*��u�Y���<��l�U�`H�x��vrF9���Sb���4;r�����f��f����X��$t��a'չk~���gݎ�3��y�dD�U�;c0��m���Q��dizc�K��3�O�����P-]ED��eX�AH�:�L���p��jԋ1�G߸P�&�C�4��!ä$�ka ͼ�*j=W�%\�їM���2���/g�d堈���,|�>�SGS�� ��45e;N�%�cpo����gm�0�"�������n�%4%/�;|_e��d�c
:V�[g�T28X��x�?fQ��=ZFu7�G� ���e��>�|��ʷƅO�L�cX�l���i)������ձ|s-�BԶ=��K��G���\�����ỿ[��Ԓ��L��~�~No6n��n����SK$�T�o]�q�sǰ�Ȍ�k0g�(z��~�_BL�]�4]@'c,��h��o�}�����V�_kr��~^0H�'�tr�pZ��o	�/�t���"5ܵH�K��VMA�>����9oVi����p���8@ƛ�z���mT�?�`��m�ռ��d�AyM���Љ��@�Bn��\��_�9�~h�(�\����u9p)��4�@�_	� ��� ��d��3,��I�93`��J,���._en�*�j����U(����5���8grpY��W=<Q�����_���W D=���t���wp }�)^UR�ҁ�ㅶ'9��I�@j���c�!��&P����#[���D8����]��' �ziV�͟��_K�@����)�`���N��c!�K�>�1��Ըw����:����P�d�C���������x�
{��;�ܭl͵9������C�Le~kX��í�Aɉ}�T�Ώ5xVH����ן
��	#D���tۇ�@A"����5	Г���5�p	����;�[���j���().ݒ�
�6���ݼ�g�������;H�`/����1������1F�pt���m��$dsBA��nyv���jp�d���!�hq�荀-��5K�{�İN��t#ɫ4�ĔYq�����CY������SbO_�)T��U����IU��U�u�93R��Ƿ�6>�e�opߣ�L.g��&M\k�# ;0  �� �ٱ_U���O"�_�c��	ϐ
R��6{� ���5�ӝy�F�Y�k���
����k^֟��+�A3+�Hr�i����!&-���0����*�����iL�;<գ�;������S*�a=M������BfW/�D
q���Ќ]���'cB�}j�t>
�ɮ����]ql�5�o�lZ!"2�g��e�������D,�a/�"$ەn�M"��6A��RЇli �W/T�LJ|��5��)�=v� �&)�	����~�ߪ�b��D��F�=.��?#��.��l�Դl��b8RX����nf@��*��:!��Mi��j��K�O��olj�y�֎��4k�o�Ӫ3H�mO�1]��<��І銢���gg-CAcih���L��g�M~ڧg���#Y_�����?,Dov�p2�I[+�Sf��� 	��V���*�B�%�ʨ�Um#����I�GNt�����(�3���SV������
-���Y�V�V>�<�@%��M�T�2]j��;�	g#����)D��L�x��@~eYo���ڂ�^/�HI��q�,F�r�¢�C���y5�9``N��1��sE7�܆l��'��ŭ�KOҢ���{�K�2�}�j�d?���Xq��6L�$�He��q���׻�1��%�Љ�K8h�$4�'O�r�ʇ�e)��-I����9�q|�t�� L:��@8�����tz{�h��b�Z0{Y3$�ܪ�G@=�4�O�k"���n��%}NɁ��_�'��a7�,r�OQ�mo�~%?��d�(�ƐA�$�Go���7�V��o,AF��a�g29ݷr�n�r�
Q�v�Wx���Xl0���^Ǭ�&X9�J�V�!��k�V�m�l깋-���}y�lD���S ���'a!Ǔ,��Hĺ�k.t%}ws7Zl�^�� h��9���j�@,���'"|�d�CYO�� s�Y(�W���~��h��t���Nmd�W� ��������̖�s�o�ߓР�*j�I��7\���^,j��,��R��9���u|�3�'�'��{�>8>#��_��4I��!w�W�����T��������pO����*9�.Co�.�� �N�U��S����	IcQ:~O�
��"�-��ӓ�~feu�x�t�bz�0�Z�үs)͸���wl�������`|������>��	w����F�.�|r< �o��?r@��s��z��Pp�;Py�Ga�ݎ��@d�N����[��`��� �=���(����<C�A��1l��Q��Q�Y���<���7
�q%Q��mk�kġ���Hu��{[9U�3��*���B�/N�0K�1	�u�y�f\`��
.Avoy�=�Wy�W�����=vy�1E�D�	M<y�&eZkѼ��Mt���Z�M�Wf�v���n�S䉒����o2�O��"_snOj���{)֙kOtϟ$��y�X��}����J	f_��)�Ph�V�,�V����-ߠ��9k�	y��b�yp,��#v�w�AC�b��h�c�]���8'w������C��]j�~8��ɍF�[t�w���j��7�n��t��ӝI�_F��^�4� [q�TT+Kbm6���E�#�����K����
"�O��kQO�~c�9�u�^u�W�R�2Yi.�	���@Ŗ��a��� �8G۶t�~)|�!uT�=�?-%�J����.3�����$w�T0E�2���|�{�e9��:� �S��6+��z�I��4�kEs��j�S%���?p�Mގ���|�AeH3�~�v.��>���d���]�G�_#v� ����"��u�?�=��4�M�[l%�-�TX`·��*��mt�aK�Ԋ��y���A�8�X�	V`�*�ȿC��Ԫ���s"��e-' �vs����m�����<�- ��������9y����8y�[0��<@dn1����4uu`��'�:)�^��(���G".�kf�{�+z��1�T�V��O
��x�g�>�Շ�F�*⫅��;J��0�>4�N��Ӭ��#()��)tHՍW�<0d�g��bN&���Ё�U9آ�Ź�uz��O�?W�І3#x��_y�N��\�y��O���Jq�襔�KO��t~h�Dn�WW�����i��
�Go�ݤ12c�uk�����5w����)�Vo�4���.j�P.�}ڇ���_k!�;�-��p�`���3���W��2x�	#}Λ�N�e�;�c}� �JE��ڕ!�j���;���Ibo���kȽ�-{>H���kGݙ�S^؞��]q��x�	*�ñ����w
�J D6,
��Y:ʆ��Q�g���$�&-.��g2*d:\��h���k1�wl2�n�H:��\.&�
����G��i�f����cL��0x�m4��$x����.K����=邷������{���J�bi橞W�6M�n���HG��ҋ-�D=�`�� _����������EUrou�(3n̓��p�8N����m��v���_,5Pkx�X��@5����#�iޅG9���[�c��_�J��
$���*��7�f�ev��������w��4�����^p48���԰o�bF�%0�?g���B8'$���*L���)�����:��Vl=0���
�C4o�~^���9��g��riBe-�6u�(����-��;Ǖ��6� �b��uQB��"�S�g�E�Va�%b.*l�g��=k��	"��(����In�)F�տ�%�3�R@QC�\g��2�h4�q�q��2`x��?.�=c�v��^���<�::�0ʞ�g<p�7��c
C�n�L����Uz����B�Gnsb��C��l�t�y=nZ� ��'h� ])��@�҅��N�!�6��b�\�󕨝����L�6���%��L%XR�Pj��\HǞ̀��ن�{�ݩ���xD����/��/�Q�^\�\�U�GG��ٷ��,'gŌЙw�+xV�)�7sQ,��JK�5\2�� +�ʋv���s���d�g+5H�)6 �v�r1�ym~��O]C�ݾ�&E�Yp �;��G5�a����}�Y�Bl��l��xR�}Uѧ�Ch_h�^��8O*~l@���
�����M����N7>�����,�y0�V�����1�3E"��q]f0&|y�r\���Ck�H%���r�r��ef͉P�̏/m|��;��_�¯�{	dS�]���}K�B� ���~V�������f������2p���!\�\�"�(�?Zg1��R�Um�Ǌq�������r�A
�l�|�<�E��*��c���)(�����"�i��5IN��xq��+��>�:XR/���JC�p�dJ�t��&s����hH�~9�Q�="��j���#N��)��Izo����.�?�s���-/Hf]�kC�)����;�����AqB�^х���M��j��+c
n!�Q�x1��:��$��=���u[����L�inr��J��i��u�C��O��Z������3�,ư�s���W�I�.է�{R�1:{l��:g$��������X�����p��1r�<��^y�jH���v�=Tm5\p���l]c�_m*����7��Ɛ�L��0m,9�;��s��.���QqX��i�%aD�E%X&� ��҈��W��B���L(i�/��H��H�qy��-�|X�J��
��H�Ѿ�^��@g��KS�Y	cfQiA�{�N6��GY�"�ס����*�$i��7�󡁁 �Ȗ'�_W��n59�
m|Vx]]�*u�x�n��Q5�H~C�����>�{�/O9D�-GuL�Q�f�q����?6D�Bq�Lɻp���F�v�B���A܁�^J(3,H@�Q�)�>5��2��+��fv����1=%Y>�g�Q��5��3��k&c������wA�W��\+\#V�zGhؗ�oG��+�^�Xq�q�ma= }�5o��9\n@Q�v4jO�����hH�y�9���8��ppVl��a�%�"���7�Qg�	@$��y܏[m�C5G�Ʊ)�c�����xV��̑T�3?�/��qr �=�.�U�*|�ٳ���H�Hs�(�\!u�f���ݻ�-1�~��2�&���kH�$��Y�0Qo��?��8�9�ȡ:W�b;1g�J�j�*eEr5Շsp�e���_'@1�S��y�?�)��3��#}��<�K�^�Jm���N����`�ꆃE�^~.?����'��B���6փ��	z!�����(2m޶,p"��y=n#[�,Ԡ��v��E����@�d��P���%f֎ug��:+);�H�� �&�zĨ#)p}iY#��b�`
�?DP���o�*N���e$-A���
�4�h��
��u�ݯ�NƼ$BbۧHFښ~6��4����T+ʒ!�,��sp#�4�7�<p��ӕϭ��<ԬJJJ�c�R̉\��N�Zx�:�� GtAI�;�	�܁S�!ܼ�N�-'��]J�Vr"�n@+�]��OӫCd��G��i7�����9��a���M��.'���/������z�����
Q���F��7����Ϭ�}�P�S�&u��鲱���B�p���>ʡp�s���u��a�|���G��aP��y�1�禘0�`�
C�v��.b9wHP�.�+�E��̉��'�3����{�y�����N2�XjH�0|�Vb,�f̤�t��%��E�E�?2��͢tS������3���t�� ��|�+����=7��%W�@���6 �\Ϛ��>8b}���k�sZ�9�Xyx�瓩�y�Ԯq")�;T9�Hg��e[ �a�`�"*�vJ=��]�N్}�ɮ_��A"z�k�AǅZ靟 �u$Ke���������_�Ѕ_N�[[]*��$3�x�w.?7pgW�c�k�j��#�g�W���-���,�4�>$��͓�ڼ*[EVt�Z��סz�򻏻%�0M�F7нk�Ge����s�1�0*8b�A�4�Kp���{�m����>���}fM���{(+n��5|"�]�l2���_#D%���:C�5���9ᔍ��hC\�����ѳ����i��0Ri�{�0���W��UZ*�m�ʩ�"B\֔�� fHW/�a!]���5�]-P�$�D|�v*���jđ-�;"(�:e�É|/�	�Y
�6��j�ߧϘy��r��d�y ��Q�V8g��yZ $V��l�Ccp��?�����Dgry��晷k�%����-��
���z�8�Ϟ������Őr�A7e`��B����3':V�R�I�XϚJ����!���9����}h�\I��	��׼!��çrT�2,Rr$P���`�1Q�D�ǵX`��Q�OB{�L���l�F�����3���a&Ċ��`8�����HF�mH��5��}�H����P�0H%���6 k��S_���Ex��1Xg��NJ������KdiQ=�'��S�aU���"q%��\sN.�6� ��yM�� #'.k�$2!��Tr��X�tflq.<R[������H9������U8I��5C`e���P�[���W�Q쫜υSe����_���80�I��*�yuV܄Xb��T`[�����Qe9F����E_��m�NC�.Lʢ �g����dځ�QY��q�y�Ɣ���5����u�����K�;�g
�'�5��l/J~�U۫��¹�Z�-��?YV�"p�%�P�I��WU�Æ`l�V�>�6ʎ����s�N�}g`D�4c��;����{7
�+�����zI�/�b2�I��@���D�g�Y{>�Z�q~��c��Z�~<��w���߅�V+�V�����i�b+y��/-�F�A�h^
)���iN�Z��ɣ�!U���c�I���a�Ώ�Z��7Y�����;������{�!&�;���#��+�D�B?wНD,���&�S
�T�UDwʎ���M�*��aX��2��S�$\��Z;�ˈm{�}e\�=1�$�/	a�"5	9��r�.��6��t����ϵJ1�d��ֹiK-Fh��+%d��FG�\XlxVHYEB    fa00    1dd0��k�<ySR�D����Ӑ-�`�R�/�K�ǙZY��T3;MIHr��e���:Ұ�)|�ś��~�b�ɰyx4|�B~��_1 ,���y �V��5����L���8�q9���K���x��f�1�r�M�yH���_ю�(��kNU{h7(�қ���+��^����h�p1Ğ�į�Fb��!���w�mU�K�k����~�D-Fd$\^����|����_.�T,�fVh��Ȝ���j�ج�u O���Ԣw�*73��^G� þ��S�E5PP��T-z���n4� ��K��t��7�O�UG�k,����F����Î]�q��$��{����4����" w�I}r��r���(�϶�#%���&�f���C0���Sp�%)l�o
L��֮�"�q��K �P���Z�S�u�\l7�3ڕ���y^*k0h��_s%Av��I����~u֭陮P�Md@�\Oweꀝ�?��hE�� Uo����]Q[F��,����Q.DYk䎲������-n�����**����R��r�e-�rn��hj���-���%�w�0�`�����c�h����Np���ir��J�_;��m�_�U�^�������?����${ȍC��ّ�%W�.@P�dP:>1iR
(@��w�'�_����)ˇ���A؀g���������y}
K�����3�o �#;m�d2��/�'�����嬃Rٚ�����i|:�����0�Q(˭�:u��,߅�:qz���4�lD�&<kj\�Ԡ���a�c�E%	^#
/��@Ƴ.ю�Lr#o3<���QlS|V4SB�k�5������wKylWSg�4�;������A|V�7���<����]��+_�b�)�l+\�E%�}�`���SZNv<�x� �F�-8ü�⭒��(�h��e��x�Q"��V���{�����`c�`�k����|�9ppt����Ò�X�F8+9�������E^����r�I�!O��[g���ӗ���=�~}�P~�%/W4px�P?� :��i�O
ut��4c:zlD�8����c�����OKy;p���U9r�d'�:�����z�Leq��d2�0VU;����ȁ�=!_��HA���Ӫ��'��R̗>Qc'�U9� ��b��9���r��h���SC�c~�"�S�3�duDS�aY2�c͜�GwX�e�k��8~m�}��.z��=����d��R]$�<�7Eh$�K��G�m`BN0fr]-��v�&���tC�}B�p�ö��"(���E�H�CU�:h��� �b�~��^�D?����m��%0������%�-q��g��l}+A0�
2޿f[���8zÜ��?���%�}AT�<��.���/���ӘNa������3�Z�pJHb(���W�n��7U�BQ��WW�m2�0��v0I����G�\���F{�k��/��0���y�i��E�� CQ�z/��(�D�~�F%��W&�IQ�:��������Z��rל0�:� g?��Ɖ��c�Nߎ	�֛�����Cx�dv� �*Ta�#y���A>s`���;���+��ǟ�O]UJE�.|�z��$0��
$e�xd�9w���^Y�&ǆ�������Qs>�Y7�%�@e�;eH�2�V�H Q��^AT)�@FGm�z0wї��7/{�FZ��݁��O�	�m(�M�n�=ӚP��GE��,�ܦ����v��y��J�Z	��ޛ���R ӝQ>��ׇ޳��5��?�eqqH�R�`�(L[�$l���NIKjH������������bg�M���fv�����W �}�;9���g-�Z�l�0����I5�b�cE��T'��s�k�;��ub�����t���j(��i�(z�aK	�H��
i�QO�@܆�d�	��j�e^z$	!6�o��Oq+�h�Ӻ��WIm]p�j�.%W�� I�	+��#���]]��i��_�40��4�'Q�t}�!RSY�� �f�V�z�*XKtWYW�|:�c���p��.\Pa�ʃD�}H�W�
ғ9)�!tV�E�j��SWO�:�<|���<S�t�*	�v��O�}�	C���Bj��a9�k��S�n����a�=���	y���`��)2>}��.��yr��Y)�c��xA�P�pk8�m~��s�F�5d���Kr0�Lؠ$j{�p_�?�a�q|��>�Z��ٔ-vѣ��z�z���-aF�d00C"vJ�	&��0�
��&N�6�����Gd�0wM��kr�E��K(�����5Y�~+)�@1�L[b��F�g����f��5�}��ΤwA��_9``# �\�l��:R�n��h���eS��X��P�@�a����䮞�5��XE��s��/��ԍ>��/��{���u��z���A��X�N��~,�!p���㓰F��C�t�e�rt%A�$�s�:��^��N_<G0/3�A!v��k����"FW�hɦ�W[07�p���ä��ajl>#�-�BNz�@��>G�?ӣDt.��@,̺�Dy^�ս/��~�7a�M���I�77vq��g���Kb� �$-EA �!p'���[�`���'� ]6:���L�v?��ƞ�uH2�h�hX$�P^#;Ɉ��m ��s�c7ٚ�����GoX3�������0��k^���S�8�� X��8x7��K�on��|��J�շ�[Q�K=0�"�����&�+���l�6�囇<F�����Ҥ�ң�cz6@g���7ٯ��D��P�M��t֙�=�2d��d���J}�r6����Z|KY໖͛���
�g������Ŏµ�ƨV=9�)i��/+�0�I�%��EkGC���-�T��aZ����ܽ$�?��f�<�0���Y�Y��k&�u�4�9龦A�41������E#��_5��Hu��!Œ>�u�0{WLR�N�=q[��=Z'�����y�5w]���Pw�W�;�������4�Dee���W#^�r;YRD��M싈?=A���@q�J��C���}_�W��}2��m~Ƃ*
���)����ۨ�E'4���l�>,��u��j�Ի�G)<�:e|�C��C|T�㕨��]Zٕ��$�����C@
�&p��(V��n�._5V�X�W��'fT�Ⳕ���k�ȿG����ֳ �82�(*k�rw�f�¯+n%�p:_n^��'t<i�ӉGG����	 ��\�aP�m��#1܌3$A=�Yw�'9E�[)�q�'rn��u[��	�d��t�C�m45`e!�|������"�4~��z���\F�"�UAry�ey5&��e)���G�婲��
���	�s�!��h����m)��z�^���]��ĺ����WX�(Z8sFg��3�o���'P��:���i�r���I2o���R��#yP��{��	�;�9*�Q�]�ݬD�f`��cj��\F�Mq�"%t����������D`t�Wg�
�8�Q��u�;��@+�P��b,��*�`l�D{dm��sꬤ�]g�/q ����M�N�^
�fIR,�8��ePs�hi��������$��c{� �d4�r��9L�Ћ�¼bKz�y�݋8`Gn�_�Pik2��{i{�6�v�T�
�i�Fc`m�m7��l�r��+<�V:]T��γ1̵�ͤr��7�j�D���Z�t�~p0&�[���Q�@@���`�V�c-�Q58>�1��{Q ?0u
������|G��#'c�$����*� hE1�w�a�V�h)��y�v��]����Q_�z�;��@�h}�]�k���.u?�2�e��R��k��`���o�cCY�ñ��ĝ{���L�+�d�Ue���ii�bZ�)"��
��0����͛GaU,���ӽ?M+4bN[���{2"s�./���t1�d�k,|aEC�,R��?`�G}���F,h$��L~�0�K�bvq�pI�ґG|��ZLΡ�����-(���6���h8	D��UDE��Q�,����'�P,8}��r马R|AS�퀖c�'�	C_~-{�_��ba��JvS6�)$��_���act�1���C�Z�*'���w8S�A}���N����4g�I��L��Z~�£��C�Z\��{���$ ��f<��]�aE݀|j���%�)�{<2ͼ*�n��U?���%�`l9A�E�Iod����Dx�ȶޗ�	'8���LǄ�[rI�������k�_�׊���E|ٲ{� ����j��Z�߱�_��\7-�
6B*!Y~#-o�7k�"��=���e��]��B���c��gVHR-��yl��z����5�hL6��s��s�J^���(t�0G�b6c:�5���Jm�U�:1J5�-�l�̸Y1|\Fk�͒��1���qH�'��KO���[���O�'I8��r��ϭ�A�W{�,��[�:G����ESN�f���_ޣT~\�_p72*����j��ݦ�딎���Z�W�c䭹 ���\�����{�-��G�P̬�hF���哒*�?��(�[�'�<bi�a�*���6�Ѹ�3�(-g����Eֱd��3@��ō�Uy?�g=���c�XS@���:���J{Z��U�賃Y���{�3��ø?v�����&�ژo�ȉ��*�l��{N��s�F�������r^��ɿ+�PJ��G���9̅<����؝��GhF�q���`L'M仼O�<za(쎈|5�OD�O�mQׇ27k�]��-ܰ�{�H�Q��ۙ�{�?��a����k�?˧����!��.�j q{��� ��5�Ȏ|���!�Hޠ�t{m���H �b>��Pn�E����ְ��G/���^��P7������N�>����Mhj������pK���V��Ɵ���v��kg�^-��C�3��7P���N��2?VOu���~�3�<~��K��n �޿���OD73��ģ�pj���nBT�Kw�m���1lޓ7�&Ѕ3
��5���b���sz���X��+x����+b.ˁ=Zx��ҭTa��_�Ժ�5�g�t%��PA3�����Em� ?3g�$�l�p%�Y�#��V	1��ZL]���\v�[��di�����¼d��N%�9��y���#���R��:kQw�l浙{]\-�*s�d�D�ȶ:$Y�.�qm���2�D�R7��k{���^h�W��Xn<��n���]��]�,�1�^QR�6W�A\<�9:U��i���y�7Q�.�|�_>VrSJ�&��+i�"I�_�.0X�@_֒�����}LZ�V�>N�hqT,�*S)p䤱�hG�+j��7�׺O�5/	�穀5v�E�>I;�r�/Z����g]�V�����@�������I~�-n3�`K��	fˑ���?֧�;q���k� �CP��y���E�n��u��������MO�[�ZN���=T����E�B詴%���jG��B���' ��N}o�a�K�w�x����~�2h�J�\��ڲ3WlxÒHB�7D�����ϴ+Y��"�h�V/���<B��{�;wr� i�⇫;��NI�hS��_�!d"0���L$��YYԒ\P��IO�ET��7���<< /��1�>�f�n��i�k#������
z�=ۼ��7H~�n�S�N`K���CS�_��ʍ��m��"7�T��#Oc�|'�TkRj4��5&�S�b,AیR�C�L4��������7��:Z(��.�&���\>d��_9�\�-R�@�`�?I/�vq�B�?��G����54�I(Z*�k�4�}�?��;�����v��1 ����+_��W�'둨S�0��0�{�O?�����Z�J�8EM����0ͣr����X�ZExf��jҦN�B^�\���i�y|����&P<(��A�Ll����4A�է�^�~�	���J��K�}���qDBR�BI�)�WX�XE��sa�7��b��9�4��*1ER$��<�%�MQ»Sv8e��ׇo:�`�ը�'enJ�� �����0�G΀��!�i���`څ����ß�#������M
~��t����H��������xB�%�W�\��Je�L8y}#o����c��Ġ�hkܱ��
P�H�v"���>�W�/��K~_ܶ��(�͵�Gۜ������ww�*a	&~d�q�r�����C5���d�JL��y^�?c])��x[hKkq��d҂�w��m~YFCtl���s�.w�tL�ڼ��;@�Ar���y?�R_0��_�όe�s��߸�ŕF�­��#`k�ql���O	����Q���so����V�ޘx��ݛG]���(��1e�n�O�č{'ŭdZ:��E����F=��@����Ѐw������E��^3v7�;��X"�����Q��i�ti����9��\^�ͱE,V�g� uޝ�������B������{�h�QB�Ml���z���9rܭw�zv����X�p�=#�d2L�6����۰���o��|㶢*�~��KcQ��~�<����];��MY�W��-��^kH���pN�	����w����T�.�%�"�53�M|���4Z��!�����Z�]���ĨI3p�:����I��1�����k��
�Mˬ���yU��%�T���!�V4"d��/rs��*����+���N�\���������v�o�y���뺃��F9�+�U�7��/돈�9F]�4Af7�Bv�G����|@�7X(-r��&��'}�#��)�zV\��y����AE�ď����B�O힊����x�\+Si��% ���U��i��������s�SՐ��V�k��򵻝#M<]=�F�)g� �a$���Cr��A>,�x�*�ܔE�+���M\o��x!iGjuN�3��`k��j��=���;]l��?Ci�m����E>�O�"s��`'��>�Y�p����(�B����0�sF;Buq���iw*���Jg�&�՛r��ۘ��}�do-�7@�u���`ò��B�엏���W'��Ke{�ԗ��³�+F�Xloa��=:��ǰ� ��s�̨@��ޮL���p�5�@����_��>�VV� ��F��7�(p�h�����;bVҸL�(*:�G��z]K�<9a�t.)�J��5Z�\*&̻�t�b|�����3��m�'������!����$ HHl6V������E'���T.	�8���+�]k���]��A��0����@p�zq߁�k��OH��o4œ��-ny&~����LSF4�ym�!��ٰ|r�15D�r�'q[��uc���D�����,�J�.H'>��[o�IU�C��j��#y�jl���`�ѣW�xЍL����W��Gh��%@��I˂5��'Ϥ�*�k�Ӯh�c�`�;w�$'�6�?�e4o*��R�	�aB��
�WĖ>���U^�N����'R����-<��
������h��~m'����Q1}�L5'*����XlxVHYEB    a74c    1290p ��Euz��� �s>��W�UgP���ݡ鲣�M��7A��~kE�+V�6�p�L�'p����/^qB����}F�ދ#��z�^3+D�����k����栶罹~݃�h�^W���9����Y���֭��椚�����zH�]j��L���������� �e�3��A>v��<lld�����^�`�bj$�K��XI��Np�ya���v����<��Kz�]��=T���ylF�I��m��Ų�a�$jW!�
O�x3*��q��$�F���n�����B�pKQ���8a�X=_ھ��RnΫoA ��'��[X�F���P"�֝B�'�v����*=���
�>�Y��1���5�,�J��-�>��m]��Z�^?�����\1/<j��,Ĝ%�AF�˸�ĸ���hN�)B#H!N����� x��?�!V��{�V)h�����+.��1�E�6OH].. � ������k����_�pXr�=7�_�m�	ֆfQ�y���B�������g(@u�9o�:&:@ y���iB���U<+�3B&`�<��a����*K��a5�����Һ�#��nP��ř�rd�^�X��7PR��~J���9�����d.4����6��Z��#1A���/M���n΄5#��h�.�/��BW�胘ۯi��U�K��6��3X��Z���@hyJ^X>܂%����N �-�~w��E�=jMRwN5{ҚS�x��Z%�$�y�������z��_>��7W���7��9#���._k�T���
Ir�N�W��̟�u@�j]��4���?˯�!6���2�����6��k°m��� '�rgs��:5-���	�،e}"3��B�|~����GV�C��Q ��g��[���%�m��'��d܂ֈH.ug]�~����IlI�$o�Y^�R(W�0�;��3��� Y�[
�x-a����U�̰^F� �_�]���� ����G�����8݊`���T$���-0���i&�3i>�]N=�GKڬ${�BBH��cо��+�,�Y<m�!SO�M*�j��YWK�	�M}y�&�8|{���Ҥ�`�X���q��BX��8z�%̪4���"�IMM�7��tJR��ϑ��Ӿ�w>g��5�t�R]a��!�V��2m����m]�l<^ )�:V���]=F|���`6����_M�"A��k�&�)h ��B	�3 ų�g���2�ݸA�}hik�'���]��`����nD��ொaihS�L��pd*=��@�|�����c�U�U���q@�xj澎��Ǟ!�� R�V�o��j{耷v�Ab��+Z����u�ѫ�\���h�M�!Kn�<T���z�4�2�q;/=&��7HJΘ۾���{2���N���}��n*�n�a�^���
�����8c�#arap�c�q����	1ϛ2[�F����������6�~+O�I�w��3�r��o,.�C�jiáv\�i )�.%���&���	��g0:3��#2�e��.��O$������8��3�uG���^t�ݵ%5��т���R�J
�5����Z�+F�\�����%9�[˽r,��`T������nxm�7�u��ΆZ�j����4�ByJ�d{��<���<[�� � AiY�G�s�0+�%*���J�&�j��a�����2\�Ѵ����o��]/6cЦ�q-˟��d��#�Il�jn��Yq�3���~���PV��U���$mj��¨�~X�RY���P����4A�,ĸ%"x�b��g�C^�z@�� 4�Lp���X}��1$���k֮�cWchjc�`�c��f|�LZ��w\B�1Zܳ6&F`7��A4&����;�����c�rQ��2��!�,0�Nr�.��/>W�n�Y�R�2�x]�B��%�8���ƻ��ОSL&��鞖�U,H��3Z>&�����߿�d2y��bs�6[�o�:`��*��38�"f�l�5�52���#oT�Ǌ`���1�.g#��H���3�xZ}]l����s.WXG9Z+��g�&"�i^]����"G��%���'XV�}Z(�+��U\/�p���/e��w4�VͱV�fc�.!�G���/	�	J�24-�T�����x,e|��;�+����5�;`����TQ?��<�9�� U(܉�,F��`���.A��h�;a%1�@A�ۖ��b���"|�5�Ե�2R�P��	,�N�vC��M\�
���TK�D�B���?�e�kC6ˣ�)�'|����BPz�α��<>C���z��N�,�2j����K�h.y�5�ԣ8�ѿ�Rnr�-N�|��QP8,���},�o���tU�c�|:�Qn�W�����P7�ͮ+`|ee�W���ǰ��>��3�p�8�qgv4lwG#Ku�*��%l�@^k�!ć� �-M�s����A�\��4�B�����p^�:�n���)�"t��eQ�4[�I����C�#RQ�n��C�$Ohw���T|}������1�Vt��X��s8C�lk�=K?=AaV�ɦ��|,��4��>�ƺ���Q������
�ɚFwQ|I�������"�S�f�w��Y�(k!������}�������%,��$���*�e����a���v��S�zx�i;�`ϸ�OW/qmR��A�M��K=M&C��T�d�#0����m/���F��?�{ˣ��.���Xtr�A_��/�5���y��8��U���_O=Itn����۽TL\y(�X���z:��"�Uu�U�~��.�䁼�!ד���N���D���h0g��hC&� 9��{#�X�w���.w��� �a�"���� ¯�8[����AW9��rj;�_k����?�"�dm���E���a���5��s��D�{�X��t#�%���G<cُ|	[�����q�9wQM�X�/p;Iç�����;�<�%UT���&�:�'�\I���wJ^��8[�&�;���s��#�v4�ɮ|e��c-DEԍ�1�ZŽh��ř�6o
��O.Q��f�9ZF���X��
��m�'���MD-*�S�A~�](��J��a�����%0��G��sՃ*v�(��B0X�Y��/��Ɨb�GM�a5�>���?���gL��X%�y
�XX]���]�+����+a�5�en�l;�n����D	��狭c�\�[lg����������]:d�}/Eƃ3k�<��� ����?�������c����fv��$�j�0�0�[T��(��s�,s�۬��i!�b�1Ȃ�F�B*��5d�yR]��B3���YU^_ܝ��g�k<,]�[׬�b�oN��.*��X���~QE�G��+�V�S���Aн`׻׳�쨃���@�&`���&H��l� dz������Q�������{m���h0ef��L��A�,U���H�v�����{��\�Ϯ��䮕�M���z+�I��g���GZ�1Kx�|�tl��~'�G/�-����7�F:~�rz��d����Gz�T�g�%�`g#ơh�Bl8c?zyuX7��Dw7�HM��'�ڽ�q��I�����a�΀��6��6��N �g�jN�����ܛ!5`�W������7
;��� ��|��j>�w��C��u��@cj8_1���)U����5֗�W�C=�,m	Fm���	oC���	럯�D���|VcO˗�
����b4m؛7�͞����au��TE��
�� �֞>F��5|�X�u��K��D\^�A$�N��퟼E���i�f1��u���g���d>�����=���ǸeƠ�K[�/؝��~� �T��dg��F��N7"8iIlp���\����!Q���a9������Ÿ2���(����Nў9}�rH���������&H~��vk�?Xpt#��ED*%����*{���ń��٨�c����m�,f��y}���,;�va1U�:2����m��ޗ˦���e k���~X!�����jL0ksH�ݏ�#OG�D��8"��=8�,ÐQ���,�p����^x_G�3@dX�c1�=����.n���7o茵�y3qy_mg=��o�0�L��}�z-�-@��,�\��Dj.巫�|}�H�*�_fД��c(n�2�'�|���_ow�~Q�W��uw�aI��@�p�]�9~:���8�[g���%��u_5=DS@T���ty�*tu��� �,d���0��/.c���Wpܰ��t{�W1+��"vȋml�'t3Ku*m�)���67M��x�m�v�d�Rig���#y�h��@w�^�^J��m3��Zk�+y3��e�����<V�]GA��[ZJ�/������ɕ�8�%�I��"�����b��\Ep-�KG�?����e$o	C_q�c'4{�i�mQ�	<�`!3;R�� ����e-�+���X��khFB����KS엇��hFu��ⶐD�U]�2��ߖ*�Q����6��ٔ��q�G���kH����W���c�����972�y �}�-�?�3��)���h�m��,wu
�
�l=�*K\����n��l�B3��N���Eʲ��4?���㲖"��M< �)�}���f	d��) ���繉Ӣ�t