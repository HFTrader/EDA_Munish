XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����=!7��n{}�iy�Mzto,�* �1b�`���)Zm?�A�ſ�bM�h6� �3��Q���9��m�¯�}���f��?d���s���I��ɻ�������q3�`6l1ţ�?�Pk�.�թO���,�};��{��D�C.�q��Rf�����5���^��Vްa�]=�2�k�|�O�g��mp|Z�y:3`��@��a��д/d���~�7#A/��˪�V$�#����↎V�O���s����8=�tfSHBE�B�v�Pl`����%�OLh�i����=�p{�o'�2��=8Ɲn0N�\T�g� � X*�.m�`:�t)�a^�C�uAਿ�� �o�	��GN�	B�,��r�G#��܌�ک�&���E���'����C.|U���!ݹ�/�Eg^zqp�6e��"�h��>�����3�a�7��j�9���������=���'<�o����:_��t�3S�m�܏���u��z��;R�?X���m9C��A�MOi�ZgOb�6(��PE�JA�J�6	�K����ߨ�x��O�@�'W䟾:�CK�b
b�b��daW��7��{���ɬ�j����t��xݳPkZ�
�鎶*`=ud#���ee;��Ű�f:=w����D��v!y+�&� r�Q����U���J�KC�G�Ns�p����@���0����dJ���2-�h`�.����po��>vX����긘�/�7K���h`�]�8��_�a�
.��eK��3�Q�;v�XlxVHYEB    162c     850IT�yd�|8�&n@�$-���Iu���Mc\Uޑ��r4yC��Ą� ���j��b���ԧ��ߙ� s9]h�k�������ε{@:��XB�o�3��u����˖��ɍp�E����1����B�l"��*����x�~_}N32�G9p�v�x�}(w��P��T�b�Xƌ,T�2[䤐]W�7����+mn��	�����E���qInJ>d��-ϸi�Zp5=��:˕�7g��Į��T�/�El�u�)��T��3"���Eyy����b�����!V�~�>��a�����ɲ�P����N2����gcƯ�����Tπ�X6wj��Մ_J򇝠Ҏ�w��BLJ�ۘ��1�|���=���9�G(�k�,$�:���K�0_'#RI� 
�#�\ϙ��9���0��ʻ��.��@�y�CPwM�a�O"o��g���s�N�|�L�u,��p�tS@B��f*�C�P4���9�}��U7��׸}8��[?�$2�3e�Ŧ����?�YM���[<U��l\`���Gf3]�#>AF�25�Xy��SH�Y>�5����2	�H��`��q��ul�8�:���{}W�jE���72��sr�x��i��֒͠�fe�X����� | �wNq��,3Pˠ)�F˸;Yp�`š�nŢ�
���g�3S����0�e�3I�j��D*H�ڿy_q��P���#��إ;����} |LVÛX,i[�ڔ��ke���ıP��c��0�}���i��N�De��K1��e�Oq�l���ka��%�"Vw�*���c�e�ƞia�qv�ۚ=�X@��R=!'���E����֑0�%����>���P'�*\�ϬyQ�j�����vK�t��f��-^�ȟ�|�&%Zǈ?�{��������v 6�U�Au4^,�tXC�S�)�ٝ��w�{.��sJy���,H,9tN���U�K6��Ά��v����X����a�E_�%������F��᱀���),���z&�l� �d,��^�
-�`p�#A���I�&����g�Z�i�<O������|��(�!9�L�����S%w���0,s���TAC�3����D���<vsD��׌�I"�o�2ɫ��J�p�p�4,���F���&S��Eӱ��"m~l�'�L�>Q�"�#�E��Lv�6A����)#BBzno�����)���}1D	g�.̻�lMx!ϭ��qn$�3�ʯ�����(?&}Z �	����s,��1��;�,�(�`���]��L@DC}�(�]��Vz2����UfUuF q����_�;��G�4<-M��x�Ђ�o�"=}�b�_4%
�-�T�	TΧ�z[:��1"��ʾb��/�4�}b���)��~y+N��"�J�9��Tf�G��.L��'��2�Q�ǳ���ܤ7�BXw[*�w��ӯ�&ז�x���[���Q��P�wY�k�Z43��=Ot{=sۘ�a���Jq����=�T���M�X ���/.��䆷�ڔa�.v����6��5����m¿���ܝ�u�����ԿLR^	_�x�[Wܶ�};�"GuT	�14)H��L�/����?����޵�Ck���l`���S[b|��M������H�r�Ϊ��NW>���oDb�Wv�����-g�k(\�.)�����N��L�'��|3��������F�0��[Ŏ����k�E�vZ�	�.N��gs?|��){;�H�Y�n�ֹ��-���N��kU�E���`bc`�*F��f��������	&�PIM_8VY�7��sS�U)�sd����������Wϔ`��˫����:��I��Z8���}����K�o���|ѕj9j<U�mq�z��G7��aRM��Z�;�
j
N�J�| ���K2�`�m��.��4���ޭ���A�}�[0�����
��%�g�l�"���H�V=�A��'�L���υ����l�c���@���A�G
���p�?���O��<%�m��}���nr�5 ��u断�WCK��|~�X�CGQ