XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!�u��c;��g,��}�����x6rp�?t��\�Xw������
b�'E���2�ͯ������r[�_��#��<{z�my˼��zĠ�Y�0ZךT�>�Mٿ��=2+��X{$�VV�ٛ��q���a�ʉ~���5��c��p,���p�H.�c�{�<G����k�$�[�6L�}ǭ+{�_���]��z��~
y��2��a�S_�/� {#*��O��?�\�[��4�<nD�I�E�nF �].=q�j!{cq��x��J�EQ��Қ�.a�]��;��r�߽r��%�[W�*tlV/�W�5�D�
 �@�[
�V+M�������5�5��t�x�A�b|CG��^,�h��1�S�����PZ!�Y���\��y�?�8@,�:��3��;������d�&���@]�&������|U��B"Sp@C�hB�����KC��[��Ae�i,6����<��[��8�����E��4iy�g�L�u@eG�On�'~ ɡ���W̼��SV��+!(�����N^��Xy(>��#��m�����uS3�F�]�'e���Ё�y��	!Ђ���� �ζ^���Y)/xI���V&A[A�]���A�/���ͱ�{ч>��Y�Tn��&;������u�a�8 H#scj��$?E� r�$Ie ГaR^�~�kz��r&1�㘳S��V��Xَ�#����Ep�X��W���Z�y!�,�;Wa6	wcu;���B�XlxVHYEB    38e2     fb0j��ONjs�tc�a>`�� �F��5fB��ZE�3��b>�qj�1,s#�
P\p��!={��C<O߷j��'Zͮ�g��'�ku���<�rO��|%�;�4VJ��`ΌPV�{���쇮'�x�?�9��� ��}rܤ��a�E_�s���~?4ߢ��E�ӷ�vJ��@BV힕1q�@�ހ��b�!(m泹��)g�2��,F��0��2�3�1:e��x	i�@
PM_��e�����_י(�m������k6u݄N�w'�7$|�S1eܽň�O�aLp/X`�C|.��V߰�Ѳ?ƭc�G�C@�)w#��_W�$��KP��'-��ޑ��>:�]`�7��ݚ{ә�������f��Ю屶MY,PN��ڹ.NC`�4���L�YY�\�L=Ej;vU�S��iͮx<6N��r|�d�̘��O�f�h�0�kJNsz���j�U���j$JH��L!���5B"�jݐE���D��z)YoT$%�6&���Z1�/u�S��*]9�p-�=c��/5��hR�~�Z�o��LI,�
�T��O���> KWQ�����󆥹��ޟJ[4��R;"������8Ԇ�P����&%BlOMݧτ��9WpC�8XϠ,��?��ٶnd��8�tv.Y[�)̱q��ʒINq�\��f������/�:9�Jx����3���<�W���Β@D��cp���kf����H ��C�H�xTEV�������fTM=�No�_5p��S�l�=�F�v�
x���x��	�Lc�Ch�,��ܶ ��xn�m9 �c40��z����LyH ���N��	�V�(#���w�)H�>�,(E<�[֮��ai��_(�R�\/��9�L�5s߉9f�1�B�Q��躁=,�tu�W��t�:DKa������͑��׀�M�� �z�+�A�Q�W�sK�aׅ3�����K���@����-�-�e�2�u��~
���7�Q�xH�?��t���� 0�/���~c���Q-�9��F�|}%S	t�� ,�Q!�bH[��)b���Az���^]��_��<��:���C�'�.6ә�����9������(�����)�9,j�6T�z`�k"�Ǐ��h������Y�L-A� 8VawD���<$�����u�;��9��BA��!"	�O6Z��C+�����n�8���VV�@���@����x�Hh����r�֖fQg��e��H�gج-ů,V���3��;��N�x�5��@�;jh�TɁ�E��1���CU`����=��,qX�~��O���� ��1��ZH�q��'��M�����x�eRAa�k?���P���9�1}�x?��;��J��=$L�Y�W�^�SJ[Y*�7k_�0�;\�����"ZV�԰*a�5����alC<�>��ezcM�x+�Ch�k�F�
�S_�dQI�Rˣl�ҟ]�iG�p���_��IKR����1���y��z���}�&P���P��;��5�v�����叏A�=��cD	�6�܌�r�y��I�޶ܹ�|��$A�������!�(�S�<�~�%�{������8��Q&ǁ~?l#Ы�w��=�ػ:d/�fѤp��VVH���!�#�Ғ B�l�9`��^���� ?���?�֝��sV�Ğ�q�@#����F�:��x����N��XLM�����e�-��lA�]�\`̖,�,��cs
Ő��^f�� �皟AiR_�d�ۂ֬oi>���Ej���E��Φ��Wl��W���;{�P�Яގ-�	B=��"�	ͻ[���}19��J�M�͝
*C��о��,�iM��x��������hV����إ ��F�7LtޗQ������~��T�7��a�	��/���E~��R%�8�Ŝ�K��[�qd.��ͼ�~3I��@a)�Ԙ�[h���/$\gƆ���^c��tSk]�ݳ����
�!�U����O]����ܭ �&K	�_u�X-yָ7(���Ki�HJi#�Yj����uӖ�1%t�I�z�C�ޱ�.a̖�V���??v��mF��0-�����Zw��Q}��a���MN�0&�<��zs������7k�0x���꿱��OW���ۊ/��i����˙;��F(�)����cO���Q�"��&���e,oM��E��I�8P�:|��-��(a� �?�)����;ΐ�)+�G���d6r(�B�sa%�z[�d�I�j6�.�J�X�r��ȳ�����s�e�	�"� �>/6!��G|�$_����
d�A��������!t��N�Mkz�iE�.��!�d)\��V�mY'�{���!��J[�f�5��.;�:i�9{����Y!�wFz��L��[�!�Yj�9wJ��!�r������Bz<�F���xe\X�6!�@	�:}8�/6���N����������^>A�㌣���Žm���_�G�M3ai��R����ꖕX�؜Z*�5&��JC�.E"�*_��/�
� �i��p#��z�_78���	���Ŵϱ�ޖ�`i�o��a�ϛ̉�$�.��V��������E��zt�wm�0{F������n92p9 T�+
�E�Њ1�8i����k��_r�zX 8���g�X��5�wӦF������;�i�8vG@+'��S%|���LY;Mb:ݍH`�,bZ��jmm������7m��B�3u�j>�D�c��`P.�+��'L9������&�2	S��#*�a�-��t��7�C8ܢ�V�(&�Ŷ�|(�|��מ��V���eWew�fS�5��>���3*�Mf�&����:*g�b�l0
X����t�Y�A��������k�3�~�;�ԃ�i��7W���ӯ�/��l�uBǧ���k�J���/�5�l%��DϬ���N8�"�pF{��$;
��[A��:��\Z�τ�eE�����ڻ���JjZB<+)���v�Ñ7��;ig#;D6N�~,������)�ɚ�P�קּ擘�R����_�A8�Y�{�zW������[��v%ѺQ_�ލ������G+'���i������]�"Q��}Av�|�h,?U�nQ~x�}�^��m(ɛA���,��>q�-3F�'^��}|�G*���+��EX�(��#�����x�����8�}I:D6�O�1��(��F.L]��p�5>9&ˏil^n�#W]�����WYS�;�8��p!8��L���EG��bdr���+�͟n��?&%a��?��\��
ID�51
#ҋ�^�5��o!6���kh�)�AA�9נ����M~f�u���2��ұ������wzi�"ٗ\�V�+�e���Q�K�Hհ��io�Zs*�� ��`�6��5	O4j#��@�!�B�~���@s橆Fa.8�K<�V�2�3Ǔ��qb�T���6�w��_��0��N$8O~�f��#G��J�H5,F�����E�c�Q��cLtp�� 뛓�	�a��ρ��#�E�U����3AbUq�٩�t��p�$Ӌ5'�)��d�#�r+�k�^�����b�ʞ��ĚY[{i:K3v�oև��k6T$aȏg���j�9u��%Pi������(����$�멞<z������u�GZ|�a�����~�{Y�䕧+i���*x�3���^�p�K?@��ebL�Xs�J�;f��Z,[��b�|fz1����Q?����Z�0��2�H�ș)�ܥ-��?�aL�iu�J�[	c{�㒮��4'��*}���0*�x��R"s��-�\h�=|8Թ��*n<_��d��r��e���g�*B���U�ͱ���k�<�n�%x�a*�q��,4�?�<��{�l3b���P�<���S[��g惜��[���d�}:����%ȡ�iÿv��q=�7��7q�	]��cm�%޲��g�Й.2��Em��