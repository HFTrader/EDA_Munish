XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0G3wl�ԡcx�Q�h1#�S����H�����|Kw_j��6�BJ��^��ʪoo28\�\��)=y�M.�'�!�d�s\PID�Æ֭!��V�����~��/��ҴZ�%Gz�A��4�C�<�';m�`"!=��+�8Af8
��zЋuƚv�"ڂu�d*�
e�	���{f
a]�4͢�3~��Rb.���]� +��4�P������7q�L� ���䥞z�<�c���-qڞ_TO��ታ��5�E� =�����ψ�F��$ڕ$�c���F�yl�&�}��nN�kDA�`L<��WyMQ�� ��X�Ǒ����ɉߧ��$��f�oj��c�7�]L,�8���_���-���#�	�ۇP� �b�§���?��J#sw�a�U��Io��h���X�BNZ�N�+�|D�&6��y���ƚ��i�
ջ�ʿ:�c�ү5��ґ"��k�e=#���"6=|*��}E��� ��Y�sr2���`�ß�ʃ�=���[�br�Ųm�f�p���cEߤ��1�����)8��]q~n�_�Q�z��Zƌ����p�7ot�S��(�U���<A��b�-p��"��ol�W�\�P�A�/��uS��3������K�2w����Fez��Q�'�\��O�����E�p�08 ���-��r�x+	A�G���J��OO�q�l	_����K潇巩�UBm^Q8��g#S���bv�>�tL͢5@(����W!���/�V(`=�ʓ� �DXlxVHYEB    fa00    1d70�����6���\����6a\3;.��Ĺq�N�r��%�t�_�;&Tǹ��w?M�]���!9�e��V)D\x�&\*+M�V�B,?Z���xW���&@U-�1��y�� Q|�t����5ڃ)�2��������E�	�p���/5�.���䦽��8�����������(<u�f��4��\�RfAM��ɳҜN�a�>�����9B^U�>�������,�R	��|�L�g�ڍq)�lX��l��Ny!b���-1���}�qX�t�%G�Ɋ���*����;�����Z�WMy����o�uJj���1S�)R���$~��K�_'6���o���xم�>�u2r�:�Bv��E�Te�Y��<�����N�\42���G���K7�$c���^j��rʹ�7�>z{[�c�ҿh�oP��/�ӮL2ِ|�GW���)��ik��w��l>�&3�O�E�0��=+��d���5������%[�dⰹ�~Y8��٥����$�����gZ���䥂�Lo�ԩ�/�Y�����T�i�ک�����@�$\�Y¸�oB�&\�RQ�_wS����h�W�l��ic��,��j�h*'�F|���a���g���ǻ��K�=��ș.�5�.0�1�n^��#"��o����>��x6���ʼ�A]`ֈv����@��.����6A��Ϫ±��J��,c��̙<*�>�rR7N�m!t����jo������4jj羆��Xkj
��lZ\(���ڗo2A��F�6�^���źC��(��X\[S?��T���}C�Mඹz�_�m���z��>�ߜ�SϚ7�duͥR�ε�\q7�'�X��7����Ud☿P����
�3��$j�f2}o��S��2����e8��O`���j$O/Sr��<v�����LH{�~��O1��M0S�o��FO3�`��.�ڵ8�������]8Т��GBm~��a�i�\K\�Q�	M�M7�U2�8�\��ɪ�n�k0ڗ2&��4p>�,�æN�s��{�x�%����ʮB��'c��0>.(�����ҪP�ϯ���t㷢�4���>h@��w��/[Jl�mw��-h�WZ�{�~i�n�Yx+ �x��k���u#�$����R�u���7gjH�b���'7�hF��@��	~�+s*��F�ۗW���}2"b��7�����������>���H-+?�l�@n�Diu�g$S�_<@�_
��.&?e!�(>'u��� w�	���3�q��W��<;g����8C]���E��Z{*t�/���
>���I\.�@4�� ����a�S�����O�|�0��V�I-9�:���"��]}�T�Y7x�%��~�D�Hz�����h�8�0,��{�����S�2M5�� ����'!�vZ��=}�=UPP�|t���tݞ���j��gNJ�qh�-D�~���g O�w�f�����V�t�O(�h�i	2A��l���u|����`�{�,�֑�Xz/B�!�w��Z�W�X�^�ӻ�$�U���|UKʡ�G����b�K1���9�c��~�;�b�H\� 1�p2�i?)˔��s-�5:g*e52F���Z��1�ŕ;�y2K�4��(�޶ß�w�y$��@'�r�6�8�WR7ּ,fթh��1��@����9�P1&&6�.U��P�`��&Ge*e��.u�!�[��$E�4:�退�� T]��L�3�l?c��mr�La�WD�F�'^k\���ح��r�C���#�_��ǒ��Rbw�9�%W9vq:7kٔewR/� Y�S_���`�������.���9���<��p_�����I≽6���<�+�~�����1�\�H��=2��9�y�?����ˎK��6���]��w&�x��J���+��`J�Ä��s-05��o+���*1 	����{HF�W�_\��3d�9s�{1�D.��_�{�4�hNK��5���7���z���\8�5;�T�u���(���bC�V��S�T���k�X��r��VL,~<F�����]R�ߧAzLZya��>*�:3g1,p �Iqb��6!X�,��:�0c�ۧ�NK�ݗ+4�;ҩ
u��(k�L�*�g��=n������@ܶ=ݔm�F�Ε	�S�M��h�*ߍ���f}�溃4w��>l���x"k">������oXj�_�k�DQ�`�W���3Fi��J�H�@|�a$++RrK��64�'g�˚y&yK����p�L)�6��ٗ��n D*��Ď)���㑢��=�"�J��N��@�F҄�T�zw�SSF�!OPC��գ>Փq�OH/ίFn��@�@E�8Q��xqJ���a8QԖr%��&�R�]A�p���~���7���g��gM���EX(AE�A�l���
�(� ������-c���#G�!IbJ����$����͟V?�($؛J��M�C��V �~@'�M��Yq��P��rff���g*򫏎*�r�������7���w��2W�����Q��Z��@w��*)���?u;����!Վ�%�z�D �rV��0Y�����9&��M^߿�+-z�Q���f�����$��@��V	~������ۯlV^���N��RH�u���2}2�L [���-�O�<c�K�����o���UR.R�!��^����C|)q��>M�cm|&+�t�6�k����� #�&ꗐ�����/pG��-;�}+E���G�}Z�^W}$
�F�F�1Fz��J�3�K�vz��K��X3��wR-+u�#�����[����T�aP���G��|�!�{�Q0�!��mǦtuzYc���C�+�;lq��bn��*9?��ZvCA�y��Çb�����F��vc�f�T�]�6��a#9���\ѝ���3�>|�w��ŏ�ͱAY��5E��e}���+���� ��BBVZ��+zd3���{�dr�.�My��u�38��y�`}c̗�s�;�FN�9�i+t%�4�V�6�i�K���Jõ�_t �T�|�,[���syh;7�^éwk�b1_ 6]0�����������H�i���8�-�Z�\��
�R�eTnM��֢c(9��`X��ך�j���U}�Y�����$X�v1:�̒F��0�0X� ?�C����Mo�|'KqNga�|�'�R���D�pQRlM����m�c.syY��a�i|���z@HGn�șw�V����&(r�6�!�,��������;7�Na?�c�Oj� ^�nk���u�N��Z����g��@�4���ZK��gt��ٝy�� ���9�
D���Aj �f:b�g���X�g֕��)K(QЬ�H7X�q����Cv)�~�[����Q$%�(�
x�&,D�m��T�r�[��a#�c��߇f�x~3sMXhq9�9kX ����-���<:96ѷ�*M�A?$��[��i��q�BD��Eh��@�.fC�`o�$j�5�-�� `������CT(���;AT����J�i���AB�_YifՌ���g4R���ps�����*�$�yÒ;6vf�C��.�kr*�D ���#6
>����.`�&��I�p�
�( �V�[�0�'�Li,NՒ���ݮ��t�L�~�%�d���]��O��E'��0]�U�?��Z%��Z�е!"�6|��x�IS�{�)��d��:��/��<̇������f��)�6G��q-�Wct��x�ֽ���4t�o����E�I��9E-��6�0���d埠IJ��FϹZ}��g ze���#��񟮬u1u����1�=�L�Gg��21Ű��>쨂@���_e��#����hK]���o���
]��n|��L�v����]���22&
���Ùr�Ѻw��)O-�p�*c��]F`c�i����`��evs�Bn�AV3,`��n����P��d�����aD�,��]��	�MDP�u��C���tf�%�/%�Щ��_dP9��x]nw��HR��0�5{@R��+���{�VD��#�cg��y`o ���Bm��L�.����`��v���7���Nƚ l�3׉n"L������?�:%��~�~ �9�mA�_��w*�k����c�u+dB�}�Dj`
J��u,��a�k
���*�|*^�p����~��>뵝Gt��G�����dz�����x+0��tu3��<���z*��_���{z=&45�Zw�ů��':$�tvod��<ț���^�M�"��bNGN�}J�>&3~l\d�Ȝ1yS�P�p��׷��9��~�ŕ^��x���9g����= i�\�#��MKZwF�9��ˣ4WG�Ǌ5��=nx��Y����K�X�kt���
���匔����		mpј;p�"��lr�m���3w�i� ���v.�@�b͂��*u�j2��;&�91Y4g"n�z"
���%�O��,�Mx;K)�<�0�P^��<����}���e��>���I�*��	 1��Tm�z-��o��[H��A
$�����y�8z��� �ˁ�ג���X�S=�����P/f�X��s@��	�P3�:�� mV���W0�@�?�%�f�Rְl΄<M���{Y|T�t��ⱊ����ksd2X.�Jd��$�U W�6K�B�Q��w[�kk�-�h4�:8��%��E_�5�cK�c��k�8����^��@b���O��T���i�p��)s��~>�il�'��hO8� &�uX�~sֆ��dB�6���e~�`���E@`�m9�����0�yZ"Y��y�<G�ռ;�!LK4E���bW�AB�?j�eZvPmROhN�J'�f(��Eu���zr/�"�)�J���Gq�����v�!���KE_Ʈm}�#�{�s�%��Ox<�;#i$Aim�	�Fb�`��7�.��0$�E�튝г�����+?�S3u㮋�0�+��N��b6� &��|��V�K��GM<\p�{Y�0D%VD�8+�~�^&�,��Y�u"�����p��I�{�;ivޅ��S��d�&�����ﴉ�D���d�J�z��U_����,	���V"O�J�{��	d��p����O-�}�����ŶE"��	JN��k�!���h~���6�����|/GE_�:)L�+�i�SL�g����s����-��$�� #�6��㈍mb$c��1���G���4��%z6�9�w��iS��L�z�} ���y�BiX�cD b�,�4�8?�i`��ƨ��^���sq�?���vG��d� ��q�wL����qK�`t�{	⟔�ߩJ'y+5
�Fbb��'⋪��i�R9l�K:�x�t�*�@F�({���:��X�,��2��j�7 �=�~�=�I��~��v͹�u�|��O������LA�d*��W	���a�f��oյ
|�M^#\�~���v��}���X${j0U�\?�EZ��!�+����^�0���D�uR?���Y���֋�AE�#2�g��W��sf�������/X[*r��{��41�x������(��[��p
x�2i
Ɋ���J���U\��n�BS=F���&���ఐ=X{p�'����G��0r�t[��(�x��*���6�B��={7�߹z���(���°Ġ=�nP�� e�����wy���/��f�X�J�)�q}�}%f"�I�~�-��/ٓ&�]�;K\�㯊���@I)���8��Ei9xe����&9�-p��t	(� *X�H�M/qx1��H!���<B�v�l�/O�`��Q�[�f�8CO!������T4��U�,��
���FС��4PJC|8�x}��R�Y��n���uL���s5V��`s�v�D�?����$�PJv�Yf�;Gr4C\E�q�p�j�T^�6�`���I)��N��,�H�W�����2�g�IiCN���~k"`�o��9Ϫx��Z�����U�����;��`dݡ�� �qbU�~H���s�e�Ii��?�7�_^*�����f�ɮz[�6l�z���I- �h���
a��n\U���O�su#Hq�U���
�4ƿh��dm�`���MI�J����7���l��0ˀ��`-��o�_@X?J�.����]�.�<�P�	q���=pu���� �ã3��ɋ ���>�*!�/>x�i��x�'>�%ox}��P��{!�F����2H�t�E�4z��%��p�v&/��P[G��v����g���# ��a�����h?u܇�sW�e�q��&�{�R�������P
(f1�w�_O�����ŢuD����0[Q#;����~3�5�Z�GT�[q>����:�Z���	�r��|y}��uˠYC��wz�?&�50�|c��&ӭ�ȠQ~sTܑS���&$�8��(}������ʐkH�"&�z58mF�c�Y�cq�@�\.D��2"}���M� ��;t�����n��Ea ���	q�n��!U� hq��
�͸�d��0A�j����E����Ӽ0m���X��j:������k�5/�w��@��qD���0y�}�7��&S��51�	3,�"��� �լ�uO�G����X�u⏂��'*�PrW�Y*��sU����<y�1H����"t����
�g{�D�ig��C�ڍ�t�8���]�ռf��E���_�k�8(v�k��_�Q7�K;��+.���1�ehY�K�&lXb���~4��{8���q:�����W��-�A�Q|1eǄ<���3T��!�p����l�������	���Wd�[0�|�����U;3Z��L��?��[z�kq��l����řK]m����+�%?�Y���O�adJ���%ι�h�Ŋ��c�{�TۇG2
�G9�+Z%����I�h���\���+�1�����fUs�V���m�v(%2�i�K&��D1ֶ��[�7�|�%�l���5̮��ՌK�G���#�c�A������ >��/�Eu+&sp�nh�>R��:�|�ؼz����o)�I�%X���,3K�}�����z�l̦�ZN����"kL*9��e�m��۹���l*���0Q��xn����Hd��3��o9n��n���KJ�#~���J�ڒ+��AS)��a��2͂����F�?���+w�������d.=�k�{I��b����14���1(U���l�Ԥ���v��p��@��\�`2���<�1]%l�����W,�dgg��z&����JP��V� ��-\<�F��<)�����0���b!2MK.����͖�!wc$���6[S�)��q��C~ۀ���޻���9�eG��M��g1I�6����a�	XNC�_�v�x�p��Tt�_��ٍ���%��XlxVHYEB    22d3     6b0R_;���}f k�@L���=v�Ę�M[+����S4���b~o/:�HE�s���ޘ@�\a'��,��~n#���:�����|������Y'0{���(kc�잂nHA�*��UAwY���������ғς���	��ώ$2���0�"]���P7t�� ����w��ݢѱJLko�[V�����˭.��~�TƘ��0��cp�Cb�����q��`�De�!���/i��NOZIq�9:�Mm��ʱ�<:؏A�եS���PS'��x�T���!�|R�@3&�]P�(�"��@��P�YY1��ܟ�v,\� A��L��~@����w�	��e��!z���E�!6�ɮ�b8�ǚ�BVv�Of0�ɉ����7�W�Ʀ��J�{:J1�xЃ�W��#��]���tP���k�q�|}ӎ����Wdv�5R�*%�'������K�>j�&I@���+>�M�,!Ug�2rA9!�a0�H!8gA�iK�
��o�	��'�ƴy�������;N���)ziA�HA�����B�;[#�Y�$|8�v�P�F����ԇh�:W�gs��r(���������DҨX�?�>��Y7Y2oU���M.A��&�ϡ��C8%���d��1�֥"��:9Uv'�ج%4R�a�t�rjvy�K���C+�@��r�[��E���O���r���\B�3��`"`"����A YԾpj�S��pX�����̵��`�&3f a_��jƇr��/��a�$0��ʏ�8�|	�*0����M���NVT��^,�y���Tm���y).:��
]]���w��m�U���]�]���&���ۑ&��a���o`�n�����$��ɋ{f�m���RLjwź4�c2�Q�!#D�RZM���֣G\2�LuRI6Z�v�/����C�a6����ƛ,���'�d!p��NJ-�7����ߧ�ad���`I�	>@�hM�<�{�2Ҝ�@��@W�~��k"���cG�<���� L����u�1�\�6�֙���G`�5�ߚi�x?f��򡦁�]h��A�*=ag1*�v�7=v;�+�V���59I;hZ;]4�A1f�~���Z�-K�$7S5�goCV���� Օ�,Ξ0{�b��(�L�\^��EKǍb������ s���k?��,bj��&8�͕w��f��qC�ݳ|��7Ҵk{T��] ��,�V�]����f�D?(�k Ԕ�n ��m���f����o_|��� Gψ^4�ɻ��*����@�A��(_��"Ўjf'�*�_�N��lqd�ڎN�`��M��E��2�F9)�����ԕ������)�
Q0�o�AIH0�C��|ꛄv�#�]c��4��׫0����iT�M����x,y�5(-�c�1���x�6����3�5Iew��!�1�{Z;��� ��'�Աt�L���3�:��|#��D�+C�3$�a-/(`0�͠y�.�k»1�x�q�M%�)��z��_5{Uw�c\�X�K��^�'�7.�9_��6q�`dV��ȋ2�3��(Q.ШқG�	P�(sa�9QS�X{���_'&��~%�]*�7a�eY"e�\[z�S,&� ��:�w�[��z\1h��"D�SՌ��:�$�����]�A��yu�<��C/Z�.j��6��jyz�f�`����=