XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b���s�g���%����"7�ٷ�,YQ4�m�mG5[����n
,eS�"_at����Hc�8��dwaX�ea	��d�-�|o��b.S%��a��׸�!����V�Xc�G�X��d~�7�m��OԳ*�(O��b���J�X���D˄4V�bhU7Ͼ�ơfl�0a���>O\h�օ}�+I�ld��[�Uye�4���%�kX��1?қ�J9?j�T�@;��\�^m�~�N��ȶ���&�mtX1� ����?��ϓ�s81r���������~Yi(�-`��`�}�\N��G	�|��@ޙ(������8�A:�Nv��2֍�=��Q��X��i�OIe)��i��A���գ�@��(�WJk�����6W�6`��,������Ţ����sy��&��j��sE���>V:ا��br@��!���G+����}��p�3����KH���#��*�S��CݳƮc~���� a�&�%�=�e����a���j�,�W���J`'z��.H�����_^��� �9҄=��<�,K\�5�=�.����߲�LV�)�d�l���y�N����~�Hj<�����^?��3#�|B�;�M��r�lC9��%��u2=�]���ే*�k�-�V�/���x�U)�����c�y�t;_���W�P��;��T"y.u6x���͵
�܉I�D�,5�)Id%��
���,j5�G��t��'�'�N�D�b&F��)�yF9{��ɗ����N�M�+�?jM��S�/~��z��ɼ���XlxVHYEB    6cf0    1960����k!���J2�,���ͯ����{(j��hS"�d0O`	C�T�����~ShPU���K�NƯ��l���
�%�
/X��T<�Ϲ�[e��״���̚�a7l���S<����|��n�o�͖�p��`���M�q��éʷ���~ �v<��������.B�4F;FV+���F;Iu�2�#{�`D ����Dh��hv��4v/_+�u��F�a`γR��%�i",_���Ք����e�ɩ�&���q�bV,8ތ��B�gu�2^�r���+�O����"oG�VoS�����$��"2�}��,���G2ҏ_g޻h��5hz�;��eN��ڭe���ӄv4I����@b���ۻ��D����!�.[!�X9��KtB#�#��>���g��fv�q�_(s�E�~f`�<2��&Yld]����_޲6���c ��j̟��F�Ծ�X� �N2����|\�Τ�`r�$���GvJ��}mq�Qj	����z�����e��r��e���d��f��$,�Ϣ�mSNT�����;X� #���W!� #OO,�&ԑV���������YS���ǜ.���À�5�|h���$�\������淩�� �@�g���=�Z]���ni�u��g뾖�������Y�N�FWe����pj������EQU;���!�9z�N$_)g�?	
�Bd 9�WC&T&��b��Hi_Î�Ps�K�@��	�����٬T�22
�7ȉ7^r�j糆�w�u�7��M�S��q� �		�Ԩ&�	4�.���r{ZP LL���Vʷ��Y���Y`N��s�X^.�A2���e�Y�$O/L��}V���h�|�5$��ӽ�:�1��V�� ����Z�|̼º-#�=X7Da�$
z紆�V)��"��[,5����!��p�Kq�ئ�+��)E^RL�.B���|?r�D��p\'TPD�S�M���<K�	�n�@�|FS�S7��4���3͈Ho1�H���'"�Z���e���gF�#��eU��%�q��b�;8�Ā�R�BP w֛�� �-�*>X�ms6����
�ɿ���Ĥ��������^�Ƒ���@�j9���H5����u.�YB�H0��phW�z����o���W��(	��&�MoMS5k����u���	��=@c8ٳ�*K�*e���q�ԍxj�'��Fnx����#��6�'�r[���}�ԎRC(�B�\��S�t[��ƫh����N�x��ڷD.V:4���rO}7�����Z��87��>fP�
n�j��#-{�#S("O"���@C�<Ԭ���z�9R+�1?`�M�m�/zlLݝY�Egs���`�[٭,i�LkX���Qwb�;i#܏㊓+��� {�����zv$8B	^MQ���߳��H�	�oMjMu���o�T�Uj*��+��.a]��/#'$cK��m02 �Lb
�)���W{��_m��������q�Y�8-dq�C�>�Ц���Qػ\��a���O�`BXj���nj��� "$8<�>�|�� 3�Mj�$:�aop'5\{�C�y�ڛ��:ty���j�?
AoZ�;��j/�g[`"��s9�	e���oVB�&�)������H�;2 ��
�xN��	8]����V�@�!;+���t!��NY�n*!��}E��"�d���n�N'1�Gg�p!?%l���ަ�q�A��-��ɛ�T�;���GwZ^��<)n�8K�F��P ��y�!��B�b���l���
��\;93�Z�-H�WR ��&��g��H����M� ��0�)�
c�4���!d��0�R� ��	�^2%n+)S����j~��hxG9�uk
pK<�\���e���~�Ǌf���Eo���[��-�Z��kkp^��� �+}�rt�[I�bx�
L\
-�V�F$�T�dՑ�_�ٞ�#�,$˙��0<7�@ 7��:�6Ȳ�[�6�ш�77s�W�~�a�؆�R�����<��5�.a��]B��'��q,�`i*���A���ڃh����S��s�k���I��K[���GO�JG!���ԢhϚ�*,A�x�N��zGo�,,�`p_�W�r	Q0�q�r;��'���o�.zL�1 �'���?~Fd�!�U�����)�B��,����Lf����ծ���7���["\���ԕ�����qzY%��tÇ�Nv �b���F��~�Xp�R�-GizQX)6��X^lUהl��Cj0?�J\@)V�հL�<M-7��9B����	����/�
��*�Ԕ2��־�58�5"�K`��B�Y���&j^�v����T�j��wb�����q{�b�Q����l<�*��ȯ1��}�g,b)�y������ io�������؀_�l���#��4t��HE�lt��!�'�O%1Ok�H��Pr�i�
Ϭd<#��&�hL-��l ǀ�1)�J��&O���έ��#�y�]e�}���A$��i�6�!��;`�{�;���������t���VSR殫���t����O �������n����tE��4(�/`n�Od�3V����c#&��U�>�Z���s�
lu<��8?�5 �<E+��nښ����j�Y{��p=K���9�j�])|� ���aoFҫ����~�����
R�Zya.����J�5���g�?��h=ïj�ÿ���κ1�	�2��tt�cL@U�dy�ZmT��U88.�Jn��_�"Qt�\�C|�S��m�%�q�Ū��m��;�Kp�oA��U�[}�D2����V���������}�l�l�("wߜ���*W�1I��K�Tjg�3�Kc	74��?�q=_�T�9�^�6�$A++�
n��8��Kીz��)�t�3\>Vl�/?R���<â���b�r6�du�ox����]�Ym��S��U`�\mݩ�تe�TO�w4��YD̪���!ɃU,[����ٚ���!���F?�=�c!~I�(�Xi!��`�u���d;�TKr|%��'i���=��T�%a�*���u��%	�ê|��|q���RRLvD�+�IOSc ����$ʬ뀠� ̮��]-�0�ToM����X����{�]5o��0�����-�}��T�cŝ��3���:{�R�},�F7틒B������*��Z,�F��m|�<V�%3�����4����-Bn�)�v՘�#I�G��'��D��T��"y�*6���j.[j��Τ��-oh��x	�����Y��R]��}���_�3M�Jch��E|h9T��m�-}���(�vB�K��R9�"�iH�̘�EZN���K_��IY����f4��th�E���
�[Q#�+0�p��hɅk��&��`�]���������Y���t$Qvc u	$��W���a��� O�;������0⺾Χ$gg��f��h���Է>nss����PXrB5��·��l��K���Rl,��d� ]z�1�A6����l�2~���'�z�'�s��>�"V��l8� �LL��sA.�R�ˊ�a�y�������B��G�;*�gNj��f�6���ͽjT���e�C/ �����R��4^a�F9G8lf�@�Wt{'\�w�O>��>ŏ�n<$�RQub0�M��k��y.p�,�|����	��k�
�|��ۀ�\��<������ތ �T��%���F�T�/0Q���w�?~�-�������m���27D\���]I��Ոd׽a�(�	��f22�����5p�f^Eu�N$O��YX*�ڪ�~h�!��F�ȃ���8��=�:�RY��q��(�	����5�Q'�>� ���i����MC�U�4	�3����,1s)oq(����^�D�Qb��^&=�5��ڊ��ѯ�/�?]辟���x�چ�4�Y��%�q��P�f�Q4����/�Z�� �,7-Y/�����0���{�R8�m-�M�|�ȫ_���>W�_�ͤ՞R0�mP��Cn�frQ�B��J��i'#(!)���NAR�%�-Z����t1?���S��7Q�Pz�%�e�:@�N��P=+R��i�T��PA?Z,j�<(�ջ�M��Q��'!k�u�X}}�T�)�q��թ�=��]�q�u�2;��;���o�!�k��`���kW�-#���I������:����+�8�H9��;hX �����7:�W����x{�Bc��Χ��B��J��M�[��,(��U�(u߅Ds��,[I�O7!�˾jS�{�pU��]G�rVN.�;I��V���`}���� ;�.*��jV-�M	��gt*9�!�f��jD�>\r=";�������t?��Jr�s�E�]���Б|n�4
i���zs����-����@������v�*����2m�(Uz�k��EB ����}�|��{��IB�_sO�&�f���.h:��1�X�	���3��£O����<�Ϣ�T�x��|yhYL-�Ʃ����q��@c,��4i��b䔨[��;㥫��qc]���_��s ��7JVb��A�����Yf��)����c�d�f���*u~�B��[�u�M���-p�+T�pI��I]���	���.J<���l����mW����L7�P���J�a2�,��@1��ru�alSa"�>5J+=�h�7���`����8�'|Z�9�:����b�p4�0Sy�z��U��4ﲟ���M�s�ƶ^���t_�Y�#��j���$2!�78o���.BjI�%ƻ�ȷ�J�Z?1�۞��������������m!�t�	��Ԧ!��fb��Cܧ�#3������N�J��*�_̬�+A���u�Ɨ��#ҋ�X����P\����:�V��MGI�\�,2����<@�-Z�	?
�f�XMj�?�{��ݚ֚9DƄ�eʹ�j07���XMS�g�h2'E���v�w<J�M�[x.5p�@���P��`a���\���H��x<�2����WO�W�]�P��\��/�^���{KO �g��]�s�NŹ�S=d��]���3 gF��3?0b��j���0��W�(�xG�����{%����V`=o�"�e9%��.�ti`���{[�6@_�Z:=�����0+��}�<��¸~��5/��������yʡD��mW�&"k���Ǐ��TV�Ǐ6ݶ���$G(���焛���m������`h��A��3��P����X��-�!XM�ni�0�"j;3ݽzQ������7@�9�:f��5����z/wi�9���H2�Ĝ���]�̒��i�H6�09��\�ӂ.�z+|��l��Tw�m�m�n�A�wUD�r�`�x��Hv0���A���}:#%������\%d�6rr�=
���QEs횡Q!��x�,t�%�����a�������	Ͳ���竁��	N�̣F��څ�O=���d'/��wz&�w���q���>&<S:f�+-�X��}[�'>1�ʝ�����Y�\{�Z��4UU�S��'��
yL;{a���a^�������[�l��Gr�'yi|�_�E�f�yz�n/�Tp�Z�g�caݝ�����h(���1u=��{���޽!G$�d1|�!���z]���Grp�8��|(!����tXh.����b�g+��y_��H`��[,���T��3��y3',���{j-���l7�WD�mQ.j!�;���z��S���%
�����buf�3�x�U)�.,*V�������3�������V2ˣ���gd�Ŵ�1w�h�{�.�PaB�ۈ�@ŧ��8�& �����rU^,�2�\�+�S^P`,�a&�j#�E�Y���Gp��zY��sn��c4>.�y��z�ӣX�\�e#�&6=��T�yT_�>�k�h=#��z	P�rS��9t3��܎1��^��(�L�$x`��bθ�gLa���l����"��@��!�%<� ���_\)3�_��{�
� �&��u���r-��H�LDxC�Oٜ��|��0�k���`��)Qj���y�vW�9��j`8��̸
d��Ɇ2f28���7�_&����.PEԭ��Ԍ�	�	YǹUX�pà�<Hv�=���h��[�Oz�5ƞl�i�V	=�i)� ���L޶���c��Z����i,V*4u���)�z���S9��)�w�~���S���2m����i6��;x�6W�����
2)�J���+���k�֡�i�&�_��D^zxA	�9�E	 ��CM@����z\k���4$,��^��/�]Rq���֔��wǥ�@�q�%
��OÒ���>�j(���.�r{,>� c�`�ى�lO��2�u���XXu` �F��LJ�Փ4w��`m	o�|�`ft羧#F�i
�4�W���