XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@v:u���ۜ��1�x(���
��:��W�0��E����T��ȧ�]���VY�&�n�`DiREW��+��j
�E��V��\���	�"�!զ�"��%$�?���Â4m�)����>R�Ӻ>-L��ˬ��jx�*X�(reh��~�� Ǭ��O��|dw�gF�S�~��#w�y��J� h�����|&�3�m��I=j5��i��	S��m����Vu�zh���qf�=����~Ǥ��bæ�zj��+.i ���ʳ��c�pN�e��g�L���:�4w�?�偕�����2�����&��g����-�(���Y\� B��h��1$�����4\�ִ�}�Zc��X�h�L� 4�KC(��atrm�ih$�3+T����Veg��x��@�|��*) t���ߠ[�Ma<Z�9����&3?�S�v�u�/z�r\L^-X�}��6&b�����S2��7f��@��C�����;�d5�)�c�4�*)��O�p�ݫx�An}��(��]�R�ࠝR�v��v��j�7lH)B��q��jt�%���퐔�a'�`W<�1UP۾���=��ک�+�����v&T�q�Y8�� s-��Y���9}�c��y爏�����2�^��]���1b꬀hr���vkn����r�T��#&'���?��[DQ�Y�*.+B��A���&JJ��d�s�=i�'տ'���y�vC[���=����3ȍ�rU�ډ4}($���!�XlxVHYEB    3504     cb0�Z��'	����I�'j��Ox��g	��5O���^h[�3�Q7��)��O'l��?����s3mM�핍`$uJ����C����U�Ԭ &�1����S�ĭO�L�E	|�[_��.����n�9(lO�6���Y0��ۗ1iu��%��`�ӷ���#��7!���e�q�v���@~��ȗ	��!�j~s��y���}:�����9�n غ�8 t��<��q������OF�\���eY�׿V����UeJ	��n�CU��wwH]�˘J�rFoD{%}����itZGw���w���9[�����C�����$�h��[=�DÂ��A�%+f��NS^	fV�L�ߴ�Kr=6���6	��繨f�:#��M9�ř቉y��E�T�F��OȎEe��(���K��T�S72�Y�%w�Yǳx�R��%o�������1�m��Lz�PP(���ն�Q��#��k_Y>a�
?���k�r�řZ~�I���#�SFɗG�Q��^��B	��=��[jI����^?~eA�[Oh����3�A�tB����9��E����ֈ��u���V?1k�t⢘�9Q�a0��5^�
�d��Z�ɏ#�lK��(DpHE���J�Xʎ�7�	R�v0�Z��rp-�C�\�;�<���zʐ��7����۱	Ӝ��[YY�ȑF�MӪR�:���' ~_6�9�V�2M�t0*��¡�C�ә��!B\�~2��[��ЊDHY�,s�R�n��)d+�T<��vs�y� (�6H��);��2���5�.�����4�\��4iI����1���-f3`w�w�`aC"ǡf	�"��W�蟳���]Y�� �<T@S`/�x����&�N�K[-3*qwie�Xj�7rA�%5HK2��p^k�u%"DG5��ܧ'MIq�x*oT���L�g���`���s�j����-`����7:�A����8X���6?Z�Y��.~��� ��e�6r��3Q�T	�=�;/���݅ M�]h�Ƭ�Oq�BO3.84�m��s��Ӝ��-)��4������ى�Ƶ$��-VsH�ۈNZx�9�T�}�l.���C-w�)yt�ieM��d @�0[�?�qja2��Zf����ӝ!�n�K�l\���L;�\��w�R�і<�]n��[��t�u_Ex��Q�9>Q|ܵ�G�u�Б�wß���
�ws5xZآ��sV>�
H�1��ޫ��fy��)����įI��D߲��.E7�]�;�3{ �f�ǭ�.���k;I~�>��)LgE�Ȱ.Lq�+�2�y�+��tB\<:ɚ����n�H��[鬎�Q��[���������:ú����̈b�R��`#姘k��H)�U;�$�P	�̴pƭ���6���B��;����TN�U��킼ࡗ�[�1�:����Trp�@�U-<�7�
N�V��C����8s�����xL���A�ӵ/%\������(�l���TA�v����<f�U�sK���-�y�D�pfU�
�q,�^�:�1�?�6��~gK�|�tP������ 
Dw'k�����<֑���<�+8�2PB�pEe���4W�,�4�|�72�<��V��0���O����O��Ђ��`t<���~��ȑiqy�fi�Ɇ���2sٿ[�:�2�����"={�f�C��ن�N���䬀x�5�`���D�1=��w��e_��V�3BƁc��#�'��dD4��|.����=�C���y��X�a�+((Aa����s��li�n�\֧�.��a�b�}_X
�����Te�:"��z�&]�M7����)L7�,��-"ʪ�$�T^�g����:���O�Ű�5K�?��Ӛ���"v>>ɮr<zL�F0��^�f�k�nb0z׬!mif��<��ꡔx��`��q�ɥ5 ��%�_�8]���J�����~s�=���^p�
6Y��75�;���s�$�g�m��0�oELp5�4��h5�-P�l�	�8+zd�3BI �Z��V���p�hc�Z�)�O���@� �*H\i4�U������^ ��a�p��
� K
$���T��j��1wĤ�_�`�Ar�F����c�ʻ� �$)'���E+��B	[Oc	���J�/����1��,�%�E��,��k����q�C�C��t��z�c8�~O60���ۧ���B��9�H�e�D�o�0��ZcW4�?5X�b�m�E�{_��bL^�i$O����;�u��ټ�溪�i�NO��!�~�H��1���6�r�'CG�JH�?�(��z�B�j:��~����J���am!����Gj�+��w	�|���w:6R����l�����F�Z '�$���c����+��#�v���`�Ǩ ����J�6�~��i��j���q$3�i���i���Z�_��l �#9;|F����T��E�rҝEVX�}��y�gA�^��4��h7Ɍ3� ��J`�?�A�����*���r���DA���B1�
5��mW�k@�4�r���po�&���FO�p�Yy-�t)��\�h�T�� ܬ�X�}�d�ym.Sd�����Iϵ�D��$$�c+Q�;�
;hQOV>�	���Y�`�SJ�);&?��,)��a�ݸ��lv�3��	������A�{Xҙd�N$�
L`�S\��^��5��x�ƅ�a�O�+4�e��e����w�h]s<^s�-���;���i�b���W�ǚ�h�����zt�Qأ��<z����%�4G}�]SmCZ<�S�+Y\ܿC�����:���*F ϸі�-y���F��i8ލ��kT{��.G�Đ��Ic���(�WiQ��iyq�(���R�q@
2����g�_��#���H�����&���k��5-
�6y&A��J�v�3���Y��><o�<QxR�-���)�mm���#$LN�$˜�}+ȅ�i��ԘZ�^��w�X��;/F�I̊a�W.Hiu��r� @��-`��`횗:$v���v��,���v�+,�u����4��A��iM.�b&g�*ǡ��U~��W4Mֹzt*�I�y���䞌�M3*����b~;m|�%[DO�
���r��x�ܧIR`R��H���yL����J2'��x-ܣ��c<��4]��A��e*�MFnj`�rat!'IE5�b	R���z�lv�o6'oE��.�/��=�D��