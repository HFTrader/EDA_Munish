XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F�Qm�}j���b$r�^�Fg�7qc8M춦j^�(���36�(���/s����<J�06���s����`���u\��]y?��z���a�#�l4 �(��"�hMUo��d���/���`Hx'rZl��/�~�
���P�C�|�-<�ɻ���d��+}5S��I�<b��g� y��y���S�����EYb��U'4�Hz�!V#��Ʀ���A&��Wǐ�pyR1Gu�P����Qh��cX��l�V"{s�K�m�7}OD-�L���i�t����D3Ҝ9Ԛ]_5�U^sH���uZ+٪L����ƳQ���0��mk��{é�;�=��7��n/7���k�W �>��+%�)Z��W1*6���ɀU9t�V��ɩm�a�)H�ЖDO)߱��@�޽�s�oO�W$�F��w��浰��:�[`��� T�W�*&z��N�n����V����G��gJPx����:j�۟_#��
䵹�%�>O+�������I�WӚ�����إ��<B����n��\�2{#u�s��lRlc�>�`���l_Kr%p:�J��,F�d-�.T�n�[<�����Ҍ��Y.��2c�雦�e�K_go"��Zgk���lvG�}='Er�$��b����za� � E�Y�j�l��\%�	�i�Y]�sʡ��T�B�Q&y[�J�4�.y˲�3@qu�c&H�b�Z|�䕗���DI|���Hn�*��ʤ6���>���Q�j~����2�XlxVHYEB    130e     7a0?F%b�s11|�4��)����܎g���M ��0�y�Q���_�+�]�X���9s�6���0y^�����t��vo������M�S��@М�b�0��c~T�jM �'�0�k�`������BX�!=�eI�dZ��l�_���]����p�c�2�3�0U�q9H������XC��,�99H��{��$y���rIک���l/�-����n�Ԟ�!�2��F�%�O)�v6hS��z�� �Z>���0l�� )?�44�IU&��@���5Qj�NF}ݏ�1��6*����l��£_�_!%cz�oWO���x�6I�~�� �L�G���S�۬��}���i@E�j�	pb����~���	`����89u��|-pDH�<��}�W��JN5>������x$8�n�}��U 腒>��</��EseV�
�o78��^��J� #�9�c�#*ԳR�Ci*�����ա�����	�01M�w쬌8QQ�1FV3M[���'�T��9�F��?���0��eK�͕�'!891�n�>Ug��?���'|�:0V�1]- P>����c��z&ě,��9���+��(�O���&O*T���;�pf��s�g���ZU��.�z�,� �d .;���
ieb�f���獢��/��C*5T��|%�"�A"��<V��s�A�&G�MQ�VR#�$�do}�ҍ��_��Ա*`����?��L̍��Qu�l:em��6���ٽ?��q6W��S��%��D�R��*�7�ޏ�, �EZ�X��j���-Ui��8P���7O CH�p��\(i��ZsJ7���8r���C�e1�h���*���������k��\��hM`�,�B&���e'a���R���0�T�|�'q/��@Fw�Q�Z�ԇ�l�v@9����1���02I�f�����2N����vۧ��J3G}�<�i�s�nɃО� d�P�. �NL�|�M�lpO�������A��m�'y�n����]i�������x_BŔ*��#��v3�AƗpY�����}��j���%\R���&��_8uxJzU��5�gއ�8D:` {�L�;G�:u"%��1 ��Y~C�h�[~����=�	UYE����n^��W7����oW�0YVdb��K��QSdm֬�ȠȮ_1<�TK��k��`��n�d�͗L�����2��k�cn��A���h�X�ocn�S-��������e�'	ޭ������EF�#E�S�4~��-�y�ۥė
6�vс�����x�0C�^C�0�x"T9���V"׸\I0�R��Y4L���n�zb�ތ���Z0��H�	{6���J�ɩg�:`�2��Д�QVl��ە�'�fR��x�w�H�@Iv��F�4��ò�v��6M#����2�ejh�Q�fOpd�G�4ꄒ���-�f�z��}���k��aײ�4�����Z.��s�o^�[&b3-�����q�M_�wu��U��~��ӗY�c��E%��$fN�����LL�I��5��b�b&#R��~��v�ۄa�Ѥ����^zG��|�L�XB���ϳq��^���b�^-I���=a�1�~l.)���� �/\�}�Gr:�O�e��H�1�Pz������U�k�F����g�U��"���g�
`ﶬX��T~d���0��u�ҧ�;F���'�~i�^�w����D���J�sq�����
��^%=KWnh����~�r阻�$�)(����f���G���3��H�sc���o#��ٲ��a�d&*���W�B�A2R�p&�s�u$B�d83���x1����*<��
G�$\M��Հ�$�U^Ii�&�E�Z�����XԵ���