XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����-�A�F��o`g��'R?�d�:c�?w��G�S��WDֈ�����ДX���q�1��]@|$G%"�'�#k{�C�T��,�8x�͛p�3"r  ���ݙ��6G�E��/�0�v�vt`��g��8�����ը%�++�ٹY5r�[F��XA䯝�o.1B��S�ZCg�O`[N|��$�46��,f��e�ajf�1?����텱b.�h�&g䥀R�\.�,k�ʱn]��9k|��a����:�7%�`���^��J�W����&���Uw��z�qduf�t��Pp��ޤ��L_UL�x9�b�j�Oh��Ƌo�#���:�S� v�٭��"�HJf��HT�eZ��� �^.���^,23X�v���D���R��Fv�+ ���(Q������R5HŋZ�0�.K\qY�(L��C��)���h�^F���ZC�Z�\�ׯj���	� �.������,[9�L����D17td��Ѫ��)��K�Z��+�N �S6�ݍ{��6X������س`����;���7�-�Эh�P $T5=T*�to��NF��&�b��%�}�`�##�0����,e�[�T#��mR��zȼ}k�>wW8�-���Ћ�ц>�!L��}vu�$���˭�6v٨��Y��&��7K�Pg!�ͭG ��n]$m��%&.5�k���L���g?Q������\V��"|�1��Ӏ��/���s6 F���	D6���.�8���;K�KXlxVHYEB    4192     dd0�dG86��2	�aoyŸ��+41Ӹ�?~͵��ϔ����\���#F�G���$�D��e�	�'R��N��tĲ� ���W�=���3���kh�H.֞
n؊����t\z�����v�8�a�Os�L����z��p'�<8ͦG����A_2Z��3��͉�P���z�T���m2L��Ѱ\���:1�E7�gk��'��R�!�o�L�*��P|���_z��	�T9�&�7�}T�Ã畅���h�����s� ��L|��~k��F��=�{KV�{H�'{q��vG��}n #���s��ʚ2}�Iz�j��{�"Z��5P��t�V#�3�(�)�I��.`��E6�#��ގlu�E'ٚ��9��=������u���_�p�Q��3���F��fJ�tt�%]��S4J|��;C<�\y�39�v�"�-���SY	͓��ex��{Bu�j�_���K��q.^T��+�QB����k��j��A��i���w��Y�Υ�薬S��*2	��I�W_M�/oa}��`��9����D9��+�߆x�<U;w�w�i]�i��0�;k�9H�G��87VaD^��O���1 �����
�E
M:��lȽrΔ&g�R$mݐ����?Y�g�����E,�}�,�S�m���*��mގ���J�lٓ�69q��2�l���fo�1�<��Jk;/QB�2��t��k�]������@i�lfm'P��3�� +	�6 �|Vu]ԏZ�����ދ��%Y�X�/P.�e��,�w�4�p�}���\_Ό˞��+䵹J*��Ff�L&A~%�F��HV(8'?���m�9Į�����K�ʠ�q�8�s���Y�,��cE��-4c0�@�]�)>��Ձ ���E�T�ߕC3�W_ �۟�6k�}�|L��}�'Ϭ����&�o�@�Oi���Y�g�z.Q�s��E�F�:|�N�MA�����nF7�i���[��ߕ(� 
3��9��-�]��oX��T58;���W	I`P��*`=:�Bm�'n�Z0��s�4b�ٓ���ր�n��0A۲H:��sX�;Yj���<��l�-صn��O���̆�Ͷ����At��B�M�v�N��,�`^�}�Ȫ������6���R���g�qu��ٺ�+I��<h^�4��Y�HA�^�Y � ��-���J�T���#�~6#]�A�kͩc�5�l�E�1�����*^,���g���� sD�?$Zw�BJ�]��dO�q��Y�/}>��
�aG#!rS��KtIۋ�!���B~<a��Af͎{�]�o�]z2�ŭ�V��(�gW�BU�Fq��P���d���8c;��f�)t���[{}.p~�)ҍ�<������?��|����͑�?����L�<�m�#�Y�π�������/@�S���wKc8ޗ�X�����o�����BDd�3�K���R����l[��5�&��}:���q�e�� j)����1-��;�
l��C���䨹D<�]�@�_7��ٯ/ۼ/VF;�6�M�$��Rx����+�u�!�4�"UJ��S65�s�e'qR*�#簸��g%bv5�sı�]���}$���RNz|8 �\�͈������N�v%-��j�?@�H�X[d�����QqWf���ݚ(�L�(S~���w�Պ.(�_�c)�>�7�L�����CL~���)���]OAaZ��8��5�+2
�h��u[�o��#���!̲�`�:���V����������F�AJ;���4a�1��5f#�m�eA���y~�H���~�z��Gi)�S��k�A�����W�{}��< l�R#݀}�o���j�]k�w�\�D���A��H�`�eX"���\���z���9u�a�2o���1�xּ=��%3	�����#쳘���@ +i(�
���>Ԓ@�m���a?�Q��x���mI/N���`<�J	x[���R2�mYjs��{�jdc�&�h�I���p6�$e���wd����6 S���e�:jl���i!�MS��c08��:[0(�JA�iֈv�.�����_��Ӷ@7�T.����fe���ⶺ4kƯa���S�����]G�g��T#��(�d�^w��)-��w�`T^VTh��0�e�]��ؗ��&��+��k��A�Җ���rj"���h�=�t�d���>���JǴA�ڊo�k�]�Fy��A�焙'�����L��@��4`w���{Kw�J��j��)J���D94s.���"���UK�H�E�&�1]�l�@1�nU� �Tz�|��YYl�����p$?_^�;��05[��d7������L��mf).�����Z���%�?�d��a��A:��<�æY����������t��<�.�����r�l�zF������p��
,u��Eu�
�><霔���v�] �'��Lk)z@��e;�=���Z�T��&���$D4� b�8�����&�ګ�_� �+˾�{�������=i��& |������s��7t p�����pQ��(2.!�o�}��,��gSv�8���5��`���m8&Ҿ`�r�C�yu!����k�x��w\���������%�]��Y��.�ڨA=7ƈ ��jW���3�Ei�z��m�l�ocpc'�V��	c܄z��^��:U���tg�[��HR5�)�#��!���p#�5J8�x�KS3xja���Z� �#w@3�eK����A��c���>`9�_\� wZ{�Ի9��@�y2!g�K���0B�%��E�����.�po�)�(I�ΐcp�U�&3,6�y�֍m�Q�:�7�e&f+�&��K���G�B�:�v�-V�cY�V��C(qW-��"�Zr:��,F��[���g��Bз)�@}F�tu��ƹOey�p��5-z�	k�;Ҳ���n�
��FD��o�����ߨ�1��Cў\�S����7� �&d��ߣ>���� �q3�*:[q\���fO]�SvW����4�7~l?d�H/�R,�?F�T��`��ƪ��(ؕ��$�@U��ݑ~j��s��Y�%���Q�:zb��7b��I�tf(�\|Ԧ��'�@a�#�0�ȓQ�:�P���k}!�+a^�1A�k�ߧ9�\�O)�3S��'�Pl\\)�fn�N���l����_e��א&��fǁHu������jj�R�W�P�(�l��E1���+!�j�9Nŵ�FGOPu�E�@hӗu��R������N�kުg��\��8~��	 ��N�mvY�T��·���ш��;��o�?զ��mi|բ��j
��t����4*�L	�^�i����h�8W��@���)`o�N�t�Y}�I�G�+͟�����2�Ժ� �hm�0�J�b[>UG<'v(�E���X��O4i^٬<H#IB���9� ȗL.��XS����s@�;fo�YI۰9��J5��p�
������%��Z޴