XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���U� �P�e�c棳LnD����QE�R�Sų~��8�R����溾�3|�+ �4�٢hsܵt.��3��~�^���n@����%I�^�se�@"�/���+6o�?�Q��q7g�_q�<�YR���L�E��W>m���a�uW����;�J�r�S$��&i&|KO�|O���ۧ'���"����&�	_�(�?�*q��6�"{�9
�����wX0�X��%���;7.���Jߦ>MmbCqDאĊ���Y����Ii�$�{��	i5�L%��,��g�G.�M��c�^-���H�ۅ���/��a󬒸�b�/�G�"R��sl�{S�N�[\���*^��Q #(���_�1� ��\Q����s&cU�*e��6���2�q��DA�B(���6�?7��m�l�Ӛ|*��W�8�PY��T��}��.�[�zme2��sw{�0i:�l�q����!D}�����{ϑ#{�翖��[����K���	�=}��}�����'3�%��)QH�����Il0�� ���6���f��������FD+B���F�F�,��ܧ՗aR܎('��[n�$�KC�nw[E��?������}��k��2�(��5�����p*I�m.Gqe�P�2h�8��]�Y	Q��5�i��%���ŋa��<�f��������1�L)��=P�ʓn�dAS1�z��T��#� ��=K����o�y�E��й��Tqɵ�Mbz�C�2�R_R����a���V�.(��XlxVHYEB    5d29    1390��8d�mWp1��ẏ6��TM�0y�|%��)�u������@"ʎ��*1YNQ�hgy�Sh�+�U��Hb��Egf�j�t��${�b�JbT1u��Ϟ#�Р�C�ׅ�r��1ց�.�mn�\f-\(>�E9�~�4��ig���"[�ކ֞��Xd���;xʞ$�p�����_���8u;A(2��X�!�~�9((y�V5�&����������70g4K���C���,�y,~�I�8�:���e���.u<��y�#TPSJ��~;�1IN$�� k����vQZ1bֺYh�a[�6���އM&��Z(k�z
M��ƍ��p7��E{��s�r2;0f�ck+h�`i3�=)E�΍��X@��5VV���};@�������E�q@��t!���cdA��%���4�?��e�)�s��Z�>/�xl�b��� K��O�T��uY�O��<[����&��+fɻφ��Bq�[���'T׃Y�Y������{����wJ�QPQ�jC�<�J*!p%����j������h�9�|=�
��Կ���8�����q�����ٷ2�����Y�j��U	vH6�0t���^^�[]槵���WT(!����J��EF�,���G\o���� �,�Z2g͌|=��<���U?Ї[V��������z� 	bx��0�
t�pB���v3�&�[��]@�
ȹR�s����?�MŻ�f�6Hк��,�m��$97b8A#�I�W�<�8�{�~ (m�!�C��1m��{)��0H.�+cu�ŘF#�P�U���-}��к�c��\�<7�M|y#շ�Ǡ�&R��w�1@R-˩5"4p���ھ��;}G����N̺��|�A�7�W�%�DݓZ6`��pܧ��5/[����xg�_�R	_QY�n
�82= �w�*Ȩ	�,K+�	�����=�����Q҂7Z��w���^wɪ��E����}��5���P;�q6��N�@f��d�;�P���yԯ��_���JW9�j�"�F��p�n�dfS�٤:#Z�K�3����DYN	r�S���,��`:���զˀ��8�~n�EF\�މw�nA�Er&� t�,���A�p�SF���:���
$�ǳ]����L�T*�1ת^���>ļ+�;v��^4�@���uyQ �J.\��1K�Hj�����bjOo*F�}�q��㴏�~G�y��L&W]��9U^۲Q��= V���|l���mvT@���U�")�&�浟��n�̺�}���LT�)Z��/��f��A��C%��O�e>��|�iK�ń�ne�Z�Lg�	���)
B/͌[A�� �:g��w����ۤHז<��-Wy�Ñ�������6�q��]��$��~��>�6��2���]b�@4V��@���S�4�a��0�������}aؿz�*�����6:��'���d��m� ].�3O�6$�Y󛒡4C�F*��:��oaN��-hu#����cpp��:!�Lu�Ի�׵o��6x�b�4��q%VF[OW�l�����x]g1�� �4'�`_�:�*���T]uw��VꏆAǊ!�/�	�RDC�qЍLo�͖�ϸ�KP�/��ElnH������S��ž!���?�~I��&\�l�)���%O����j<�8��]��)zj��?^6�]z-����QQ���0������n	�#Yo�2���>��-��Qlh�ǜ�Z�������mJE
�ޗ�Re�[�ʷ�sLuߎUra+�<$�V0�zZ��m��e��@{2�N�gm��O���%��^�B���˘���`k���ԇ�
-�q�w�%���֌j�n�u�i�
�]��L�-�X.�}ٖ\Z��ˊێ�z��V@`xs��ύ�4�Ā��v2ܺ�Xzl��VN��˖私~������>6HJw�8pΓ�Jb/7AB&E��=��7��6���Y1����r[�g���X��>�O���J��h/�)�jw��K��F�M�43�oՒo�iV���[��nG3�q[G*��9���_)^�i�l���	��x�|�G�����\K�k�����0�[.���4��f2�J*(�ܕ����gn��js�h̪k*�{�{�3恢���h�Ҋ� ���P԰�!��5[u�u#r _�ue"��X�\9o�����1B%mhX�c������)�߬���jTM�ݩ�Q�Ur�/TK�Bz;G7�a�Z,G�k���mJϿ��8��
�o^BgK�3��	�C���>x+�*,o߼|�����XV����
�aN��\s�:U�E�(�f�d�;������R�2S������yE��:�+���~�|Q�R7�W�V,�ʭ��rX
���M�+4R&_�0�A���л�F��M�!�\���tąBg�y�H���=����`.�Y}�ak%o��479gUd�^�
P����&�⥓q	8Cr([�D>�O%�DE�-܍=w����07c�K�>�L��Qf�1��7?\aY����~�&� ���WJ{���r��BE�HCTϯ���]_a�|pY5G=�E���/��K�ϊ���P�j�r�n,7.�}RpT
W4<Ԥ4�o����gC���ޤ�'����-An��^��=�Kn�P�{%�;5c�sƼ<�1��QR�?P�@ˇ�!vu�ϲ�ɔ�-TQ5��-�/�\t��t��<揉 ��D$�o�
N"�w�9u��	���Go��
n�2ڕ9F�b`�P6��?��(�l����� ��sLY:�,6���T�E�S�6�Z&`~k&��#�6}���,*0!�8�"m��(��?c�Y#'��&-V��(�Sa��]�2ᏺ�?Q���_� x�9����M��%��H��M~��<�ũ6�piRd����:�2C�"
��h9�]R|��֝D��=p�N�(֬���ß�74�����Cvs����]npp�tF�J)�`ہ�R&�֧��$դ�@�[�r_%0�� Va���}?\ȋ��*���A����h7[J�h;�����gJ��������~J�%L��N�V{�z��ͽXjy�,�n�0�	�"��i�a;��]�O.���h�@���?ԏ�T�'�+�+�?��4�8Ta�^{�29�g-e�}E5f��cA?�X ?�:*�m��{ U����gS���@/�yR���Z��9����!C�!�$^2�&]��Z�_��}L���{5�Y�0~ϻ�S�ќ���%��¿��Oi��H}b���mӪ�q�t����������P�|D	)��-hf��۩m�A�B�o{lڽc�].O�s�PК~� ���n�����9�i���ɾo̾�@Q����`�ZK$$Q�	��9@�c��ħ�-˨H����o�ϲ��wh�\�;\��[�T�_p���R��-��wS0&v,/��R@�� ,vb7�B���B�ՅMI]/����c%�Ҟ~���nG�� κY6�
��y	0�o��$T��s��z�z2�t�Ƭ�J����6c
r�@�7�.ݜ�x^M�����o�]t�5����`�6Dlok�u�:�WsY�����7b#Q��Șk�}H�����`���޵����D±�Ot����R�'�2���耤AEi1�����U����YG�r��ݟf�2��邼j'C�ml*J@K'��/J����+�P��"o\��`���J�-��Cp�A��-Jޕ��!<���r,��-J41k����!�Y��Fv���S:!h��N���h�eM�uA3�v=rd\��b��y�h#���pӝ��ӥ���VC�?hǍ��hi �Q�8,?��.d �ϒ�����������+�`a��Pܒ����t�;P�t��!��t��	�x�g^Ad\e�O��+�+�&!��j+�����ÅaL����(I�.(��Y,ob�a��=�YR������|۵D�t�,�"9J�p�����?�,��nF�ug��:�G�j�yW�_<٭s�qR�(H3�j�9��1���\V�y����������H�ܗ���ߜ���F�ӖQ��o�Қ6]�gmv���H �`TG�$w�x]`����1 ��G#`��\B��Մ{�G�0�ܰ ��x���n�]@�l�)f�	�  &kv=@j����)��jf�]�o~KR_��*gIr�}�1TˇP�>s�-(ѲbQ�n�C�{p-�1�����p�*��	ݾpu�L������Ed��k��R5*�i0���C��T}CD�'����_(3���\қ)�s��#~R��GKk3�/�R �Jԧ*��͔S-(.V/]�S=������e!B��`�����x�{��U}z_��2�,(�+�N�6_:1�4�s����(�V 1ݲ���B+��E���M��wBԧ/�\�b��L�uZ6�/�S�{m//�Q$�~fL�o��ƍG�sXw'�^c�O�(78*�2�`���5�j��\�]��X�ŉ��r�AǽC�>�@	Y^�D��?���pgݺ'O�8rjz�"��K��lS}���`�!�-ź�˓WQ;�,�V�(���  ���V��K��^ӛ�j�)h\\�.ʐ�GƑ�LH���j�fhDHO��V�A{d��K���#1�4A"o}���j@���jk��+[�|U�-�zS�3��"�r�#H.�&'�e�� ni�1�p��� fK��d3A�k����gA��&{�����	��!��9ݮ���HrT�Q�?�����o�펱�EDŪ�K6ڶ���;�
;��5����Ti��v����P�a�Dҭ�!#����\
s�ި� ��L2�透�mj���*7iz"�2�	ެ5S�wM��\��]N��\==U��8\�qg>t�ڄC��_�����ļ��^�0��s��r4C��7z�
|-�b;W|G.]Y������j.��I�]�D