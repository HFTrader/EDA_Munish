XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1]�b`�Q4B�]����ѣ��1�r��M��
�q�Ps�x)�{p�V����5�y,!�߮L��vrɩ�F*�F��A?hB��U���<Ub~*>~�3"Q����7���XU��h�,�����c��<3����{���~���BM�ד@��f���LkF� .��A�PPV��a�L�/�� ���a�l��MX��f_Q�rȤ��&� Y�M�#���WB���XeD������R�A �u�PB��S���\e��?�,W�ٹ�w�J��YXL��2ಓţ�C������ǂ�(㾵c]�Z�6�I���,	~�a?�kI��B�/�>��#d�֭�.A'½3d�닅�qDk�\������;XS��`�z�����6�<�K�n>
���/=I魢곶*��_S��ȥhr��u�n�ۖK8ܐ��*�?$�WU�Ȟ{gT������.e�����g��֕Y'�\\�HFʘ�"�������7�'b�܌¯�����zi��,*�l_8t��1�	6����-T��[�OX�G�~Uy����S���t6l������>o55��O��-�Ϧ�4�!��N�oM��'�z!�*���"�a���25A�,�K^�	���̄�� Gn�����j�}��B���MEl���Sd=1(�v<�P�����r���Fk�G ӣؖ���3���;�R2Q��"kPO�'����$:�6g��L�O��i\p�������qbJ�XlxVHYEB    2cfc     c80�:�:-� ���A�n�\�Y��yk	#�c>�7�S`�#�o~sxx�8��/ˍ����t�fv�����Z�S-֜n�`�/��E�+����J�s���y(��9��cįzU����S�ɼQ���]la?R]�l��iz�X9->J�49㽟������󓐡��H���xf|������O��7�>��,����|�@�@��=�;�@٫�77do@�
�H�m��Z��~�\�D���F�ȧ��h�q���!���X-[M�;�0+�bʋ�]d	Jf�=9�t8VŁ�%��Ü����8��JeQ��Hu,��=���\�=�CΤQ'�Ѣa\-�,*9��
�ouA���/�X.ڴ֮P�4�wCk�6y��Xړ��B�}��z�f�˥���o�;�Z��D��j̻�����ɦ*d��,���:,j�'���wHD��7��սV����&�3R%ґ�7���`���|�H����	���6�|�0����h��.�%6��%�}!�z��޼U�W�v_�`��g��_�?�F.͕07����^���\������W�5�˴�96�ǎ	R4�D�����W$s��&e���Q�8�N&K|�i7{��k�պ,�D�m�+��󽪕e-�'�N�v�?�U��3A൙�O���/9��:V�Q��:����G����M�Wx�#�z3J�j��<8r���QoN�_�@��Y��h[,Á{�׮b��г�;��1:�P��*{��5��������y|맵�\`����-�g�DILNM���v$k�	�x�����Ί��Ҭ`�����aG�p��%��a��O����y���_D)R/��3��i�p.S��CN���ul�R���:z���P���ĳ`U��(�]A!�V������w����o�F�y\��!Xw� F�ƪЯFj5�[���"���JτC�o&}�V*��_�X��9��r�4h9�����8�8�z@�lQ=�w��x{�_ͲB#+��·�R�!]�Z�������k��	%�Ր���Rt�{Az�q�#�y$��垩��7��؝�;VU��)LX�x��eCx���hs��N"��X�0Yr�:-%�4&�O�1�TC������އ
v6�{�SGt��H\�p@"*b�R�{~���qh$+���U{G��	ߌz��PZ���]�fB�wV��˶��FIs5��������Xj��^r�ɏ��q:I�iЋ�<h�9g*��L&T���*>8���?����FP`4<W����]k�ܙ~��Z����P9B��%�g��C5��5��X�وa�a1μR������\9)u
E�l��l��{z=_e�^����1�%'�C�0�lZ�9(�ޒ��^GY�%���Է݊���V8PR�s!.���'11[X���[
�o����jL�(.��L���Q�^�����.@�Gl30��8
7��� t(�"��u��2?F%����{��4�բXO�(�y�`I!��n\a�{!�W++�Y���>9�G|^Z�a����ƴƉ���Z�~d
���#o�-�ck~"��$=��ĝ�>��gdW8x�N��9��� ���E����nP7�1O�M�Ld���η�s��o��[��~�����7���%�=F-d���5\	���}�O%P����h�svzְ��_	�&*��B��� �6X<�ͷ�&ޖ�YP�
�:�Aw���v7�6�i���p���d�CO��i�7� "��&g�|��	ae���a�����^�r��V����?	��$���Ͼ�7W^�X_���B3H�х���iM�ZF,��E���KGڕ�f*� w�*�����w���ȩ~b!1�c"�܅��G���ODBGHm��|8w��ʚ��3����q/�&�7��b�9�w�2=�(�T�W�"�ި��h;�?�7�����C�o_�ǌrP�%K�i�p��7j���*����j�!��M�g��r�0���qT��8i���7a ������Z�R�k�$���i~q���c�=V��j E�~zS���YJ�[��w��r�����gy�5�N)���(�,Tg��*�+�x�r~'�T��;�p�+�S8���U��!�Ix�;I�~(>�xʣ��zB�ZԐ�0{��S��"h��ui z�x>��%��m�ٍ.{�u�J�/i�P�����$䯿��s�$�z�L�8}�c���`=Q��1��>Κ٧�,��l[ʃ(��VØ��̱/���E0�6y��J��>![J��Ca:��37����;j�˪���q9�+�/�)�e~j��Ɯ�%�Z���*j-�1֮�<,Ƥk��>"���9G�s�'�Ʊ�r�yQ�YL-�I0�����S��7�(���G�{�2]<��'WƊ}Xu�>�H&ޞ�=�n�8@_ZA:z5�,fB<t�<�S,��/U�'��*ß	m!���nF����G�ߝ0��2�.��v����L�Fٯ�V:nC�oH�۹(4*��1�Ē��wt�|�f2���}��w�r��ۃD�0k��i��@�|4�\@#NQ�3h�g�ؑA���,�A��~g�;��m�-�5a�̈́�|�Iĕ*=�ա�T'�VwS��my,�Ƅ%�O"O���	�_�2~��C� �Y��h��\:�Λ�SK���� �w���$ӷZj/D�UIs��[*Z���\�|j��]�Q	2Ȋ�}�G�c�( 6�f�H$%���	��[����]��/�l�(��#zo��uVDCM1���)��ڀ��%��4a�VX��3�^�ɅKNPMh������^�̉aC<���Wq̹�ȹx���Ž���N3wJ��~��Oh(�-��_U�3���b������r����8��⳯�SsvٟcUy4&O�3KL��(.�i,Q'�)�g�U����7����B���f����`�c���	=9O�?�5Q��b�!��Y�;y��<<�kwx�c��qo��9�tb �F���T�:e�2V1����3��(�9	�T�f���w!p�v�� 3����q��^Y���a�� ��h�6�ۏ[
�&4�p|(��VA�P ��#�������/�M}V���+�i��0*�