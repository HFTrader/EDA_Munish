XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��sII��Q��^�o
��#o���|�c�h��'F���s�&k��]�]�'+� n"o�,򯲝i��[[�1A�Tck=^C�j
Gl�����)�s�!ruBY���&���V,���I]�^��8=�K܊�zt��.Q� �ڸ���Xކ�?�߆���o�3�cLs�.P�:ad�1,wC=E�-��#jh6����^�G�f3��G��H�LzJ	=l%|Qв�]S��~&~���w#�-�#ޙ'K�� ��~J��`c{��������@!�G�c>��4p�\�Z9�7C�`��tQQQ�'ٰ"o�'�f���M��4�����s�`���+����9��<�߁����眆�ސ����.�@��
M�>ȉ@��� `B�����{��լ`a($�֣s{ڋ4�%އ�����v��wv'�e�	;�p�\G����t	Y���,�݈KX}��I.�l1.Y��L��,Ҁ�w��^u
���V�U��Y��1��競fF���|��t�<����*�hd�$�镦�j�+��w)������!�[f/����H�=����Bg��\d����$6����-�#T�}�|`槷�r��X�j-���"3���Vd7�m�54�<��*D��K	Z|�v�x"|֡�>Б�9�4�〾 4�����H�@��A���b.U�9����9@q��n����:�I�|WՊZ�%)"�T���6���]t�-��ml�G�XlxVHYEB    fa00    2520�FKZ��{9�`�t�S��!WL��+��-����$�^�,�5� �q�~_��$U���0�A=�_ɼ���R[Z��g	dT�f��TrYĪ����x�T;�fx9����v"�_W8��кDf5�->�~a���T�q��T2xi���BT1J�՗gCO奮�yw�r��g�!*�F��+�'���rO�&� J|�%��Ԛ��ݽݴ
i��m��Ár����+1����?��'Ԑ�{��v�b��(V�1U������@�2�s�@�����i�h��/��]���p��]H�y��ޒhpn���IM�w��̾�ԝ��F���"�!M�$�(*�#]b���7,���e�\և�g�K����.�Q�J]f�P�#�|KΟk��X���DP"�Y�"; �_�.q!���s��Z�P��z����06U@�����;�g�ޠ�Nac���,x{��(�E)U�&s��x��ᘽ��9"n���Xؑ+e��O�R,�?���7t��ʆ"��������
ć������kR���WEk�hѼl�-�YCT����)���{��Awɫ�u�����cS��<�w�|+�p�[Hz��=��K0Ou&fz����;�� n�!�������h̝��Jh��ɽ����y���_�p���f���qBUc�@���ĸCo(��T���1��FY��*����l�ش�����1܊�Q��gV���U�
��D��
2S�8,pS�� �{��-��e����#k��;����\�t�au���D�����tx�$ya"�l<���ћ��wG�=�-;�~K �an:K+�ata?&�1�k��r���1O���� �/��O�ɼ�Tw�6�M]��P�;|d�Z_�t&�	�~�Hy��^5��P;B�<�7B����K�ߴldw۸ơ�o���-�aL�fS���J�]�!�>	�vtM�lIL^�=�t^:)�hSN��I�-�1<)��>^fX���C�{R�U���%�H��m���"��D^+u��ݯ�"���3�K-��H�u�:����g���vh�\%t7K �� 0F����L�?y�[��*�n�khqH|Ƒ����fWޚ����S�]���Ҝo�̻�D���;6
�C��z��H�|����W������,�G��93�G�tp>����d��նg�z�t�c�x��}(x˺�*v 5wC�xc����x$"e^������`����x��͇8OQ,pM���p8��ښm��h��*�
�,V��Ϩ�n��UH/S�i_J�P�Fe1��*��7	;���{�&�5��݂K���\�\a�o� :-}�?na�?��R?3�Ȕ)��J����g���FEȘ���c��t��	����T|f�ȇ���S9uރ�y�p����`M�=g���F0���ja�O�;��%��c�O��=�]�B�ޣԱ.p��@�:$��`@�R��$R�V3�5�HX�|H���lRD�L�ja~x´ן� ���Z]+3e��L��^�?����(�͓�n��\�'�Rh��
.oV�8���Q��~�,#���B|A�rE�I��Q{c�d�q�,�=��p$7�k�Afz���in'G��&�����	L:3>��ߡIG�n�G,�aY�l4�!���C��N�tQ�v���+4�Hd���]<�]4��K�|�y�>���q�,��M�2G���9ɼ�2�=�(�.�d4�_��y��Gk�\�O���G����7�!����v����S��&��ݟu-��HH-��*�6`\���TX�N�y��V�E�:*?E�i����qh��&�Ͼڮbp$�W8�F��ꖺ�6n,pw�8[S��M����|Z �Ɉ�)�	w;H,�I u�r9�wu�2nMkX<f�Zr���8E2߅����	O(�h�~���S�-�e�s̎F/���U��G~�+���/8�b�]~Z� �^�쌓&�r`,��+m��£�����P8���c�F�����=+�/�D��Jp��/���d�pC0�!]�ߣy43R>��S��噟:&L��c
�(ϧ r��@W��I�E�]�֏��Խe{d����.U�~Z��H�����wf�5~�=7���0�P�n `E��M�� �qO�� ����|�0`���;N�<p��*}l�A�Tk�I<3�»���'���jzg��/�|�.�T�f/6��IX�'�9�A�`k��ܺ?H�<o�0M���7�v��u��t��s����7�۵���I� Q���_Nƺ�9\��n��Dx�,��|�-�Fj� �Řbv�.��	�n�,/ţ��J���W8KM�~|���#Y�����P7��`�z]K�;���S�<�T�0Z�)r�\�4��&�'�h�z&	���iݾ� ��M]�y%P��*K�jo#��� u��|��Im!r<=�)����C��ĳυ'�O�֢s�d���CG� 1-��s�U�إ�p��\ŨK%VE}�5g��8P��/z�H�&!�#�i�ha�&�5+d�WZ&خ�:��_�)����/�ի��(�0,�?��թѝ���]BH9�wI��Q��=��Є���MNo��r#����P�Wo�0��"�����+L�E$r3�8�Ff>x���CL�:�6�qje�w��(�ϱC��9p��o�����E�vlZL�M\��P��-��g��ܫ5Mq���5b��J��
m������wy���(~Z?�Uw����G���(S�K���Cf]u�@d6\T���tpOeR*-c����RlPZF�W	ɕ Ie�Fr(q*����/PYנ�;�$h��U�M����6���jX	�|���z��e}��j�ET���u�j0,�?�@mc�~��n~4����@��hz+�Ŵ��������R������8�S����MU��Lms�_�I�L���g��CVKsk��PHj�җ��Y7~ºqf݄G��������d��:���μ�����51c�m �$U��B�q��r���	�Ʀ�Jm��C	�T��&0Hl�������S9���p��(D;�vx����r��T˷)%�'(�ʼ����_����*�,�R"�oI�%^�>�}݉�H�wt;�z"6.>� u>�N*��m�xC9� V^�y��Մ�Z�ؿ�@WB�@��l�ѿf{��,�����d<�Bp	H:S?��_л��b�Oa;�V�ԛ��z�������U7�{`�ǥ9�$B|����+!�J[-=������,^E��C�;�߆�{�Zڽ}'wK���5[�zC�	����.�Gi�Z��sf�BA��6W���F���*�|��(��=�Q��"#�7�r�'l�!+�����=՘c^AU�嫛��#�=�wV�}�>F�� SV�{MX:�
Ѭ7)��ׁ�ŉK��Œ��A�u�}�Oƿ�����5_�E/��g��c�2�@b�t.��>��ʴÐ1pf	���s��g�ԝ����n�^��<(���m"&)�g��J�4���z�>N>�u�d9�����>�dO)��e:w_�OX��5^�ɳ���L�=�@ؘ4nb��xf��{���kBu�fvĸ�<���6��������r��4g1b$4V^�u䋂�]Y8�!l��K����!*I9��V�����{�.��X��t��K�9��/��k���rV�v/�i�b�:1��[\� 6Xl��M_��s���]]��6]_�dڬs�n�(7�q������r8��r�ʙ�Ƕ�e�Fs����#�̓]����Ʒ@!n�HX��f��\��ȁ���s>H�I���}�ux��S�������A�P�/Jʣa�5}�MX��S����_�����}��ga��c���. 2OUl4u�8n�W#�,a�%��#�]�.�Gt����_�Zz��wy��n\?[�._#>TT�\
�O?X7����[,wP�I�?9i���A{z��]�evk'lOQ\�އy_Y�>�7�*�����v1_!S�����6�H�ѐ-1�8�3��5���	�e*C|ro�I,R��B�����I=e�٭�n�D��ؾ F]�y`�Mp�إE���&����0J����V��%T �)���iQ�؋���C	��4�O�l���ٻ���v����T��)s���( ����Tp����)T]:�A��h +�ɋ&�Č��/\\T��#��'��Eߵ��e1#�F����0���Tv�i�� �n�� ����LC��dcIȅP����	��K�ά�F���hX}�ϊ��u)������J~�u�v�
���"��T�D�+����e"�c�٦���\�=R�W�r���.�^�%�r`�TO�5��ڣ�Gߚ�H-�X�A؇�9<$uZ|~@�=�;�b�a�)��?F�䄙����a�C��]OWJa�e�zF\�< �c��S޸���r��&����K�ʩ�G�0M���Q8�(	�4�B�4^i< '����.~�F�r��M����	��'�չ  �k��F�m��޿ud�8w�����b
(�xu�Sj�yq�C[{�o��P���)�A���#��)�Y�Asj��L
�[!��p��O�35�~ӿY�C�HM��XΣ���"�������DS�}�H���Ŏ!�b	�4 ޗz�����QQ��Eӯ.8���m��6(�"�͈�?���v���] ��b��.�D5���bCOm
v^�ט�+_�>KZN�%�Yc� <e��z��Јy�D1e���T�~TH�aWQ?�h7��G�n������� n��^j�v���ntq�7�_$~!$*8���ӭ�}(d�׀��#d �Ga`��g�Ӟ�0(4������"q����_Y�j�xT�7�ʤ�|�.��aYC�0���q��Xn�*Sg<�z�������m��{�W����� �L�f�a!���F��Wy���c�R�dvzvl�:as��7�[��W.@��l��4^P8�UɃ��w��j���#����`�r>�|�`�u; �e��Z!|�<5�ǔ��a��Dޥ�gr_��de���9b_�}��܏�#0_+Z��y�1��{gN�b���S�/ﺪ?�r\���R.�7*<��y��w^����D� �L��gJVw�(Ɩ����ߙ�c�����r��M��߰��`@��f�F��i�|.� �*]���"��ڑ�J�X����
Jh�{�4�����h߄��,�%�޳�(�k��8��x��4�t�Ϳ^�D��hh|?����ǹ<�(HRN�W�t��NCi
�P�Z����t�V��"����M�,Nx?@��Nlg��>T�i��a}}^P;��e�Qڔ޳/;��=���d�� )��D;��M����OZ�B��xȭ6g�8IK��Ƃk[���׺6C���@4�*Z����n,*caN���F8,a��m|��i=57YAt�e*����z��/�ޫ��C���@q]G�6�X����a����`zq�v��m\>@�oʹ;�g竖��^M�q���%��Z��u��Җ��(���^�_3o�'���<��*cǵy�aR�N?�bV����D��Rp��Y�i
���YoE#9�2���tpx����)dQY �4{�|(M��3���@J>+"�G�;;�m�KK ÔM��n5,.�8}��xk���G�$� A������7}��$Zq�G@I75SݝX�|�X�5��e��f!�*�_>�kzU��ݦDͧ�~��x�[8����Q{6Z��$(�e����GL0�3D��p�N/$C�m��	`��3P� W��E`��9;�x�dH;#��򹡵C��Ǐ%k�����6C�ڋ��D��T��r�ߪqlS���MƦ739�J�$q'h�	-�X����I�T��cd*#��J��}��7�aL�,��3d���cQW���9��$��P/Op��M%8E�1�9%sW�C9�n��v��'s���:ca�C���3d<a�W���}���U��[_|_9������aZ8#��\|n%A�帩kC\��#�:�no3�(q�E`������(= T�&��ܭ`����I�ԎF�\�A��d)��B@O�e
6����֝��+�f�_��0_x�u���K߻Q#��Qy��Fx-.||���'��
D��!�Z��X�5JR�}u�;Dg�q��!��8o Pڿ�9#.��Y���o��a�#5V >�G��t�*Xn+�l �m "�c$���M�^s�OK��N�[�m:{��J�P�6d�w�n�y�6Q��G���5�Q���Z<�0K��@�3~ȇ�	p}
�Ұ����`���ؼ� }a�
[ɺ䦍��q̘1�A�����޾��9̃n��O�2忍�aܖ-��~GO��������eNy�%�Ѷq��z��j�o��H+�r(g�&��#W�̫�f��\0̙(�(�v?u�y�n�Y��D�r�@jӪ
��Y�5>�-�`~P�L�HO����5��<]��+��&�2��X�y�,����3Ue�B&�X��ǪJ��G���K��{��yIZ]���6/E4&�/&g�?���}��FE�d�{��c��dL�e��/i���ˋxS`� �����7hMˍ��\no}���FW���<��֎D�fAlk�%Өˢb��{?5�l�xy�{���	oE�D6K�2͑���q���7�e.�ؾ�D�Ѐ�����F�}����^#�����7S��||f�.��0��}�N%�b���¿� c�Iq�:��S<KL�5�CщTB�`*~��+�Ϯ��l'w%;M!c1���c4	�O�>d��J2��~�mv�"{۰O��(�j@�8!�#@���g���<FχXsC�"����y��`s��*-�F�X���Z��OUo-����hLR��$W�#G]�4r?�y�:�NK����s�[��,a�<�B�L��.TE׃xq�w�w�܁-Q驻j�1�!�ԵP=^p�K/kF�l/������p&������J��"E�5�N���pebn��ƥ$����DPyJk*a^=�E�� 0��)�l�cL�VIk+33v=�`"�#ks�p�N��{`G_ڍ��;�h�#���Ш �Xl�`6�����������V�D�RO:[` a}Y��K�pz��h������I�!��Ң���c���FםH>���,�N�MG���E�8��m�:��ޣ}R��ˈj�;+"�DΏ���wDAh+���:��K�XY8����!�?p��Awmϑ�֏�����v"	RU��(�E��O2�/'7���ܝ���p���&��(�Z�;��o^���n��X��9kS��D��Q@Yw�����(�éT��zfc*����]^�H��D�ñ
ux�p`zsI���)�7E���|��x-�t��P���:��q-�G�Z�����_#$c}J�H=���1��;� �絶�]$ށbbN�V�ld
~菛���Dr�Z�n����'�	�c�U��C��M���A��)1����m����e]M���&�	��s�,���n��4P� ������l��6���4�|6}���	.�w���|����2��A`�Ӻ:c�1Ɵ��	��Y�w�eo�$���|�.풟�7���D�$_a��w	��s%M��{5X�M��	'��0��%�#`�#��D�7d���Cӱ�a�Z���e�s"״��&�Լ2�v�!����qIeW�!��!�/U<�����([W�%�)���,��uА��^�w���
	�e���������{hD�HN�1���!�ހ�����g���S��k�:��&��2��"���*��8QHܴ��f����y�m�����Z،ּ�}��Y�=��+�>�7����/"ݷ�*�~��������ğS�K8��3�{W3�^�/c�{-��Ҥ�6��>�^�$��~��O�
�J��,��5)�^(Z )�䳢�I3��;�c�Y��]�?׫Df�h聄z���/(�NXg�M���%Y�(鞓A��[J���D�	d&/T��������:�Q��hh��.�l�>�h6b�?����G�^U�'��ڕ��٥qpԢ}gx���p�-,`�J��Y���t���6GH`�͗[0�,�DP�R�����]��� K[�d�B�1��N`z�X�L������w�Z��
a�#��`�}o{���_qơ��J�F^��2�z,��𧻓��0�9^=�36?lb���b���iz��7�l�f4|��EE%uUR%�� ���+��?���j]VN4!=;�[��!�-x��n��;�C?ʉ�l���|�ϧՍ横_�hS(q�2���i�k��e��J��q���p�ͬrX����Ԟ�mL�=��3�6����
:�V�6��ĨOu�/%���(�{�*��׉ӯ�0�
a�,n���8�>)&bIi㏪��b��dz�����8\�hgl�����?���9�����t\e�H�m���}�����3x�q�OX�s�g��ϋm��|�L���.�S��q��J���Բc����W�_1�!!��L��f�'���b��L|.���,5�"\�f�!5����/}��!� ��+���|>�����p!U�wBВ83�C;/xQFspq��iM��P�)S�xU^����&]�=w�$\�<�Z�����XU��D�a�>w2"y�"���Wh�|��'"����ӐJR��`�� ��1.���|�R���r��q :�˃��B�3t綔!^I��XM��Nk����7{��p��?h��[��T��A���_���h��.�[{�X����":�F�Wy�#_V�W�$��%�Y��p�v�g�؎jm��w�%S�1��EP��$�)�����򠳺0?���[cߑY܍��k�ﳱ�\Wx`f}�R;��:�ߔ
2-�'������z����wm�f��=�y ke��oz� �g�:������L�S~�K��<t�����z�Q�l�r��B��D�̉�!��VSo%�Wɵ�>%�3��q?wM\�#��9���/�,�����?a��v���)�X/k Ɲ�9FD~*sKM�0Q�\OEkѲd�i��'��3<Ox,7���i��e�-v�WH��+G+�<�T���R�ag���0"�%������^	l�n��	3�\��RS=9q7 V,��U�NG4V���~w��7
������'A-īF"�Y%�����Gs,�i�q{�,���׆�1���_#�4������l����~��?<N1���oo�Q�"��)��y�R��4q�xm�kq4<U5�}U�)|��D�&v�{Ɲ!L�#���L�+�EXlxVHYEB    fa00    13e0*��K��X��r�6m�3$R�бE�����5�PÆ{,Qݦ�e�=ѓ�ޭزO��H%���0�Ե�_[s���p��z�>�[�;�D�1���E�JeCɌ��#{����c�kt�cW6��"�g(��#N��!xl�D1���a�� O(c�A{���������2S�y�zI�����r了�#P~���&H�ߗ�s�B7��-�������L�c7VԆ���@��}�٩]�_L��K׵�<�����h��FzczBn����g��F�����n�14���|w�wਛi�7��s��2J.�yz饌n�<2�xUЯi�s�ey���zn��\K��u��g����t5������͂�������O��U�i�Z�->����p�~���q����W +��A�,�d�H��F*-�Y�8�ze�����%8hI���H�$fT)��H������_e�����zi�h���E�7ι(����� lձ�\r̯V�o2r ��,5蟪̯o��c��և���!���`��#���J?7�cѬ�m�z���M�����>h=��Nu��AW��зͦ����d�'?f���vc��- �F�+�02ɪ���ŏ�5�-�V�������� �:�����atd�?�GX�� ��R�Jy������� J 1��İ ����Ctq�k�g+S�R�Z�}�H�&bK������u`g�mGs�DP�Q����=z��Jf�h�YJ���5�QW!yT��]v�k!Gy2�j=5�{�?�4x�g���E�C�3��
����E<3u��AI�P93z�=k���s��">h�Me)��( 㦍K�̵n�3�8������3g��	�T_��jG��h�B�%�p�7y����^ ��	| ����l"�ǳ��k)t��>�������0����i����{��靡��ɆS<sk�?�~R��0�&��@���&o��>_X��KPXa� �
̕���q�/���#a��<�����ъJ����l3�ɣ�׬Z�ܿ��|��RM����������I{���!�k�e����o�l��.x��fo�[���4}�|�f�Q:*�<���� �p`zM;e����nD)0�����*�@�
_.W�4�)hT�H�x��$�p~6	e��۳n��nS!*�l�TAFD~�n���)r�9�d�خ=4�%�((��D7�i���Z��ePTn�-��gʱ�ܿ��Qu7�Ci?����%��Z`�TE�kҝ͒fY����Y+�s>T�9�I��xS�Ge�r�#G��5�k%�C�9��q��j��e:�V���񔞡d:e��@99�.L�k[���M���xD�sP�ݗ����Qx�*K�w�h�PY���J��衍&�����ɐ/���Mt[�>�.6;��gT��^O���{���v����	T�EG�b�̺�UZ&HL�8��@��\��T�����Ad����p���H�Z�sǚ���(�ˎ�I��yh}��x."K�J�?���/I�إgg]���,}�<�i�&���97���r��ѡd&Xϟ[�?'�b@�@�i�u=G�kɣ$�L�,�xY�:�s�=X=%�p���?Dd픹6 �����"}o�w�DH{�fn�h���I�3�`c`���h��8���-V2��A�G��@�("[,?d��齈��`;'�̿lֻ�kNF���	���a)gD�C&��q��4}0����G�>j�7�(=����̈�>^vZ����k��B�m£�;�w�Z�i�M��+e�cݢ���u��������C�+�=��DO6	c�Zt��Ï�=���t�%*�|,� &���g�O����W���R����U���L�U��z�^2U�#U����ݷQ�J��6Yy��@i��J%�;�C$�E5�Ǘ�� ���G@'��>i �A>2�y@����(&��wOޥ�Wt`1	���rE��4(C6���ӑN�e�����n�5_�@�wj��O����)��W��BuxlaO,�?�xW���D�_�A�%-�G��� B���颞�ti���VJv�'g�}y|��G�9�p�^��CR�tI{."�!I�3��`�q�eP��k���lYb��|��*�ET�XPNY�J8SJh���x�DdgA�����&������YsB� nb�/w
r3�!��O3|%;8��O����'}�$�5�iy���������d1#��;��������dN�$�A��B���!Gm�|_�ݖτ�eh���$��ws|K�p�A����x�ܲ��U���?�E�҇)�@__��4 J%��;�>$�f�����1*сqԋf��?G�ɐ��30�ݒ��c)����ʑ��}�|X��It.�!�l��۾0�D�o|��ڟ3�1�k;"�>�mL5�y���e���B.���UU���:��V�Gwș�^�Oɼ՗�͗�>Ɖ2)��HO}W�@{|`�M4�8ʬ8v��2��L�*U_�.�O�]8�?B�F�K�qو��2�T��S�nΙA�V�_���H�C���O[��]#�Nh���g��	)�Q���,U�5K�Gr�:_ ��ɀjVs���=2#��JK򶔈�8x�����a���+�*�U���o]��eI|�煫w)�$���w�Q�'6Ƣ�h���J��*�z/
�m��FY�P���_�J�*D��C�{ ��(Qv��h3�-yߎ�a�������}*�c ���2ݔ�Ǉeiv�{��h� wIm�=�St6��u7��>MlL����5C�h�E��ZY���Tw�}E��sT�i�e�������^u���?����-5�k\U�N(b�=�o�ZK�ӓ��K�as-����P��:FS��v�>2�&�R��$��>3�d�MY��I�R��\t��P��L��~}OH������F���Z��̈��}m���=F$��WT���v�DI\�`��a�5��Τ?"�&m�3�{-�X\��i�BɾZ��J���q&�с�Go搜�]��=[�MT�E�����8E�E�y73��H�XtLΪM�p��ྻ���8x���`l��$i���l�?�Ӂ�+.��X�,��u�!j�e�*9�R}�˸����t�/�<KDO"4��u�tg���O>)�31AKV�B��vܕ��X;�9� ���|��I�j�
\;�t��a�fY����
s	�������2�y
/.W+�9׊w k�e��]�j�Cis��橒�	����Q�$A�3�����|,w���>?���s2�M��j>_���\41=Ǳ!�4#�@J���K�8������Z��q2Q
��z�����s|�+��h�b�W�LÖ~�Q�;�M}J��{���L�tZ>����s�Q�%�"e���wڹ�!%�\֗{�����X�ΰ��X�FUH�*�v|�Zx�^������ٽ��D�����}t[ote	w�gM	(�(��3U����sN�Փ�6=Z��Dg���:x�)���o��5#D�f���<p[���}G��Ï=���p��:�n�24�0oU��"Q�V|�v�}"6=]�ԃ��/�d�C�K!�r�h��%t~�~��zt�u���$<�6��Rg"���r��:��z��J3˽��+e�=��S�e4�T�-�Y��O�vEm�jB�To �[C�m�҇9���`M�?yM��O#Z?_�׳yp�����:l&i��`�eP�Q(W��þu9Th^��"�4Qq����Wf��Z�0�,��+�!6nɡ���ZC�o��[�S�"��N!(�,i++���CfF�/��cc��S�Χ*������֡��g�	n�G�`[I`8p��e�~ۚ �l���u���� ]���C��4�7�R2��T���4�!�����:�3��SV��D�W�"�dodf�BX"
}&eᇐ�b�0��j��ykO���.d7���V�^��y�֞��О�_�}�W���}�8�"{�����Z�4�y̵���g���Ӗ�+{�#`'�Ϗ��4w�g�I�2�8���un^���m�R��4�M����R��:�8B &�fS���� ��𼆬���JI]�[Bi���?�ׁ۷�	؀���$�KR:�vW�i��;��&d����έ&�3<�>�?�}3�.j����w��i/� ���I���G����[�#8��ݴ����m�EH�O�Y�4:�KɆ���E-�'� �\P�2�S*�}o}����K��D�x��,��i�FP�t���ė[XF�s<q7�V{ה���;�N���h�Y�`B�y������#�c�c!s��|�h�ۋxi����û�����րѠ�j����ue��XQV��c��h����a�A@Ԗ��	@Ŝ�>!ƏE�f�$�Τ�)@�X�Śzr4�H�+��X�⋚��~����[Y�����L�1Ω%|��q��Hq|�L�z&��0��B�Ix��#ܖ�Z���#.�6�8�����R�\��"W��~`���.�C�����C�����H"*`�_�f��x�G��Pu�V�J���m�z-Ӫ��>N�:����<��z���n�a�i�(�z��2`��}�1ˆ_L!&�ߕ�%���f��hv�����y\�����󢾠^�_�0V�&��7�/��r죗/�T�`��E�|k�ؔu��+5�v\@{'�he½w�_1�"~d���^*`d�M�o�G�R�`�A����)��mA���h���4��Q!��]<3¾������9����J���AG� �������u�
�Q��I4����R#��!�m~p���fe�h���lg~�M$��̌�x}����<(�z$l�$�V쪮K��ن ��p/V���l/ꆜV}�PM�%��SF��		M1�.����)�{��ԯ��߀�19��3�����b!z;����<��g��"Ol5o����(,���՛G�U���6�#Z�d���u�|K\7��=��y<���6�W�"�����|�	�!�y�XlxVHYEB    fa00    1780�~��ȹ�0�4ȭ�v�<+�/��i��g'�1[�{-l���F��2	E�k9�u��u�Q�'S�|�a��3���r��#f��ˠ�/�7�;^��Q�G����+S
�c/�e]�����I��@�o8���,�p�I��^$!q�����lϗ�3�ۛ�i_d{P"C�=�"���y�vp=e����`j���ڭr�>19	��:rC����r����"=��OV2�����R�o�ރ���� �,���,ۦ�J��D_N
�t�#��"��ޠ܀;\eV�@쏵�F
x,}�&�2Cln��z�OSH�tD�g�̈́����ƹ>�h�����8�K/�q\$�=�����$ˀ�n�%]2]�O�n�8�7�A�VOézO �
���DD�P�]*��$�nNy(�u�:mk����.Q4��INV/��v��=�s�#�Be���	+R^]tY�"�Om �����?�L*E�gqqq?��1S���j.�d-�����|G<~�1���;�&\'����\���%/��V;��1rx��6�Y�Fs�,P�!�u���y�Eg���v�P���R���wa�J��+�Hީ�Qޑ��6I�hV�v��V���4��݋�ӵ��"�!0N�y� ��X��n�����ǀ=�͐���(Ż(EY������`q�$�]��]M��3A/_��:�BY��y5��LTE�!Q!7X����ÔcVV
uoj�/xgR�w���C%j�|_��M)9�g2��|����$H?+�ENzq�H:��'�rb})a���uB�}�qM`�7�\���-XX�k`����*S.fRo���_�!g� ��]?���2����T�YF Y�;�@Q&�#����y�Vi�V��BAa��x���@`JCC^���DXy�N�:Y�a�۩,ߩA����E�����m�8�T,tn����z���R%qf�K���3t���k,����VQ¾�y������蝂�x�+��4��d�|�՚�}'�ࢠQ���_vl.�p��[J�hIO����V9��1�zx�9��^E\�4^�E7!����O�d�/�'��Љ�a�o^h�]���M�՞^��I$���t�e��$5Et�Qֱ4
c=����ZxtCrP֟�)y�-�1Okb�R'�P+"�R��p$]�gh2�g�h�� \�����"����v����k�t⯋�oλm oatǋN��\s�KBѮz����p�܃ƀW�pK�7�F	*�6�Hd��?��}RO]��Ҭ���y�:ᘐH����l�@Bj{�hA����AtdQ澋�0% �ɍU���,��)x�P�"��;b=f�ϣ�C4��ٲ�4�O�w�G�=_m�Ϥ��0H�(J�T;
(�@H]eSJ>P�HyY��0�2L���V����i�p��(�ϖ}�i;�~�𕱈`
��T�(�
���5j�f�y�����L���m�'no[���'��۠�Y�9x����'�#B��!g;����"�F�� s)Eb9�:إ>N�r?��,2nm0�?8�%ǆ�O�l�0�j�g$����;����W+����g
��=�WU��;�G�M��[��oV��w�	J�~VFxW�a�K��q<%|oVA �����٫U�Yk8���� 6��t���JKǶ��Հ��:yJ��P��m"�;"�C�����.T,>mV�r|As׵�5{��)w�>�a��%��&"֖�&4�)kU�5�U�tat����C��	��v�
�{��l�G�UX+О�T�:~��v��z�X盺t.\2�\H�An�4=W���{l-\|P������"�V�6�� '�"�_�o�����}��V���(i5����u����k�m�ouQ�m��C?�����ٲAO:� ���<@�<���l�4%=�(�I��an̘����[���@O�}z��%42XV���݀�x�/Iҟ��=���ŃR
�(i�\��U;>��F[�e�n�1o �pw�^���L/��K5�1������]�� ��gG��`.�����>,ʑtѳ7�d��vI����Z!]�},����6}����uZ���:ͧU�h~������>q��>\�x��Z�d���×3:�7�K�v�"	��h90���v�2�.�]���4�U���m�j�ڛ��t���c؇nǰ�|���M��}����r�Ha>^�����1~�*r��"�ݡ�!ci��T�V
hLf��%b�����u �S��̨��G��u��6%0��02��WFgUS+���zv���L^�?�;��E�!�Jo��@��u��f�������Z}m t�Q�,_�T!$x�g���P<��w 	ۘ�?���}� ��3Q��7�j��mX�<=u�-�w�d�w,a	1Sl�}�g��$�<�Y�-6�yɫ_�1p�yL� �W6bq���J�����S0w� �����cs���БFoD죑T0��6�zT�?(K[��;e>3�}���u,|���*��V�j�"�Ye�H<�����v>/^=k\��Bj��%����U�S��Wz^(Ý�)��'�n�͜��"����������c��֩z�����;�p#k~��"
Ǟ)���I�����묓:��L=
�HB҉"���A�X/�|�a���+��~�������H%J���@�^���ft�È�m�d�R���SZ؛w��@Ф9
p�h�a��Hƿ�g�8�h��*������.A6���(,� 7�������bF6u>ź�I��+�S;{~�-U�Cך�@��86P��~��k_%��&��� ��o�K��D
�d6�Ij+��61�5�e��[�y}�ҁ9(��Ux�!v%�J(D(5k3��W�#���O�K$�C1(�ܿ�'�O�A�ALP��Z�x+%�a��	QùK�x�1P(ո����*ĶU���>��eL�^n;��D��N�0�)�u	m�Sa�����)���a���^�m��؞�	M��H��-�!$�5��}o'��s�pO �Ez?-CA�r��4�W?=��݊��#	�{�h#r�g�����R<��R��-���J38���3b�Rʔ��`���zZ�i���d���	�u6{��T�^oc�V��Eq�&#�Dm�=����f��\��1�V�qm�!��8q`bO�����}��Mu@�hZ!i��㢘����{��?�I�;�V�f���4�͐o|6��(�}q`ѤA���w�w���Q�[�á� ��t-�3cۆ&��!&|)��T�z7�-�5QB�H�5@�Xu���O¶�q䱌�3*���&��������of��`��	�wgR�!�ϟzP&6u|��ʸ+����'gN�g�^�ؕvg����	����r���-����P�x���?A���U]�C'P�
Syb 3��Q��ME�=)a]+�ɰ���`�O&@,3cD��F"ZT2���6��w`�7��T^� �M��2�����vQ�U=�Iw�1l����;��p��싟%K{�����}���I'ǘ)��V���C8%w��!��oMP-T����Bx�CdO�i	�u+�d3�<~��x굃u��دU�̹2+
 �ְ@�Hi3VFG�1?�/��1���_�����_�nB��Hcyx?��`)�pCc�e$� !�J��+8j�v�.G�e��t���?*�(ND�Y�w��'+��(�⢀BH`zC��:�03yݏ[�/2ܙL�G�"��4(��m� We�I�	%�+A�2~�
$���w�uՁ<��И�7x�]��>�xyW�k	j$~s��~��\�]C�N@��b�=�Q��-�޸�KCJ�f�\�)� �#���i�(�֭���mU!h�̗Q��ٜ��c�q�O1Ke(R��-�O{B9�.˨F�;�F}�oJbցu���b���8[�����Ë� ��H>�?�H�%��F��w�y� |���yTT#Ne�������T#�����C�Ku@i��j+6�� 6W/��i�@��Li/Z�E\��n(�Yjme���Mr�#27��u����0���K[���u���-_W���h�.ّ��US��&/B�L�sB��������V ����ɝwlUɈeh����T|����۵�� ��n0�n��L��c38�UǛ++�.�ϼ��$�?�`����b�q����?����% ����
ܴ2v��bN�jg�+PvV��e����@s��]����!p�Q��_Y���	���[%��t$�,��H�u[�{JxZ���@ �:i�vsmSs�QX�eC�k�n{`ђ�OF�a^*A-�V� �%N�?_R�FU���j���}Hx2��\x!7F�����u;gk��;Ap]�ߣ��Z�>Gi9�X����;����.`j\Dy6����g�6J���Gxg�4Z��œ��}^�%�A���J��Mp?�J���NxCd&�d�l�hߟ��$#dG{�}��G�_�b�8��ʯ!K�q��eO-˗; :Ms݈K�{�E����n1���tS%��7��lE���?¤Kh��t>�@㵻H�W�q�Ǵl����3��4�a�p�5�ˡ�Sz@����ł��Y����,��u�U�S๡�X�@���bM��l�ډ�57�UcL� VÏ����F(�N�%	�*���S���5Ҩ*�U�s�s�=����5�\���\���'�ц�'f��M�#����#U�)�1xs�ME���~F
�VB���-�[~���U�d��+��#�m�`=ua`T�c��z.�FR�j�`� c2�wS�JVU6*����Q�wI5��oe��]x%吔�ӥ%���JV{��K�g�@{D$O<B[�ˀ2��:u��N=��t_���(���[d���}�<?4n|���J̘�]�8k�4)!Y��Ǚ��/&n�=��vO���"�y|b憎�j��b���4���W�� �D.����=9M����ǈ@!�����q��5ZT�N�B�q��ׇ��=��	8��cV�vC�Md�̜tLZ�H����yR��X���keŏ�P�)GkD.���2�`���g���,v�H�>�i˲=F"�pӗ�D�^�@��_�p���
]/ryx�VAi�i�b�(�Pq:pߓ?e�r��ϴ7_Ma�/=�ʫ�z�����ݑ>a�a�����v�f�H�=Ryu��K}V����a��;�E���)�ݝ��y�y�#�&)�7Q���6���v�^RdJ2��� f�JaQ>	�Mh�,X�X:�Z���E!�}a>��P��P����$�qg�@7Y�0�c�\�r:mo<�[/�^�AZ����{�(ق叄�ոx,YnK �k�U���I�jy���z�q�^쥝
��M�C�	�k氾���f3����z~�i-q'�B^����	M���j-�л_K�!Cg�Ʌ�̚�U)���P ��(��slνb�h o�/b��G�y���Z�b�ڢ� ICYj�cnq�n���Q����Ȩ1�8��C��B�g���l^���jWu����'	��Y,�p[G�ê��E[�}֬C'� 8�]�ң�M*Y���JΤJᎅ���ٳMҔߠ{� ��Z�έ�ڋ����L�c��y������0��r�S��%�;?�J�l�!x���ՙ��+�/�߀�1��.��ML��@�:�c����W'�	��y�L�Y��1������$Hb��kf>+�p�Y�[ ~Ƥ� �i�t�n�!)8�s��鲋�\4�������P/SF�m����SD�册���>R�S���{�X-��Yjpd>B��4蓭���z��N��v� �D0!��,����m7Y�ǡˎ�ׅ��f�r�DyU7��\f��(|&q?ՏY������T,a�uQz=��>��*���F�&ѡ,�+y/2XlxVHYEB    fa00    18a0��1yH��f���].��b�,��g�}=wc�[��|�D����l��֯颪;.�U�F �Zl�`�!�������S���x�'r��7 y�[�헅0B�����l�BD^6�M�t��7L)�+�;�^��1*@����w��Q�x��&2��4`Ϊu�q�fx_S/.�Pkb�ò�ƙ��ɡ5������*-eɯ�B(!�y��D�Q ����Ji�~��?,��cw �c�.AH"�N����Hl3r!���X�AC~I���������Q�P���$)m�J�u_�D��Ğ]$�~�1]�$h:���8[��E|���U��� Q�	tuX�U�Z��Ω}b�]�p��+R@d��?�ViW��8nP���T( _�4���X��4^5jsDCļ�J�M��L�t\�3ÀG&���L|"F��N�I}���`ą�1�(6c_׍�H�?�zۅ9�d'd*�c��,"���D}�k�9��8��� &�?W7�MC=-&@h�y��\�l)�c_�r���iW�աS�&��7�Ķ�H����&���e8��Y���6��U�Ķ��gy憲�Z� g"�|�5!S;e?��N��?w�#�2��(N�C烢X}��-��=�}ҰqRD�NHW���4B>�$z�(y92��R<O�-�����
P�NJ(>k5��&�E�l2$g��Au"���\�֩�p߽�j�#2�ߵ��h�1N� �B��X�ѧ��d 8p�H����!�n���*cR�����v�}Q�n�G㙭�FR|���z4쵅�WҞ���w���r�M	��� �#K=�G��f��Ծ�W���am�3B�!��xgb��۵$w��g���C�&����['�W����9�8M�G֫�d'p1����B�E�m-��瞁����c5�>d<md��W�v1���?���� �'ŷJb  ���OA�cŮ�SʺxzcZ�0G_@��@�ܶ�:����X6�� �h�S5�$q�}iߗ�JX�\!M���7@0�#ƕ���bbL��XKh�6��Pw��/�e���'	��UO{}�˕���$�Ʌ��$���hO��M�"�ʄR��<rFU&�Ҿb�w���7c.hܲ&��$R��VJRl�ϴE�Y˪�\8��÷�*x��{���V����c"2�R	E�ش�[�m����ö��a�@���ەX��N0��f�a��� ��QG��l��4�>����˿�C�����W��w]�d���o_в�O�����M2"��Ϋ^���`p���~�Đi�Z�4�!�;��w����fs�������i1�R�9��x/�~Y�7�}����|��RD"ʈLj;��j��v��sF]��ތ2��Բ6����Ja�:�_����u�k/��q�r�:٦VTF�B���j�H:L����-%����� �'���.$��6��.�gd;������UMG�A��@ut8%z����cɢ�0���:�+�#΃5q�����snw1�l>���'R̗é��g��7���]��� �v��_4��quK�{��w���{N*F�T��� ����1X0�:�]��@� |��Q<hk����5�t_��vQ����w�������r�$�}�b\H��
g�IƲ�vg�l�ro����bʜPԌY�em���xX ����8��H��?��D�I)�D<G����П|���B,�s'���k&�E�4)��:kN�p��."?��n5��i��KVJ�?O.����I�%��X4�Z��ۃ]m�,�Ф� ڄ��
��֍��/8Y>.��V&�?�k�R�wh���L�UN�^	��ݹ�%�6\���!�!�"B��]ڹm�d��Uʗ�+V��>����}[O�/=��R�M��diZ	���a����0\o���Ռ���7�ť�6��P�+�1�vȧ11�gK���ĸ�pY�<�x=6R�҈j��1��נӧ�;m��tu����m��yr�c�"R,]��6��p�ZL�V�fE���h���5��:�v����+�����x����TE�LKjG�St�GX���eRm��ӆ�$�H^v�>�9��"��U��+���}Y/M�q7@.�au��}jO��`���8!K��╱H�sO�ׅ�/�.�G)���#}X�x��Y�p�bd����E؈��h�V�v��OT��>��<,�wM��|ѧ�D�������F�M������  +���
���އ;fӇ�'��|&��UN�:^�^a�n0dZ1���{ ��Ӟ{{�*�\�a�;���VEV�M!B��Mx�;�$�l�(Og��8?�8�bq�*�}f���'������ć0�i�����!�O�ˤ�M��,���-�d�Nƴ��d�_�J���=F�8l�ǜ�1�d�O�#I�|W�=ޫ[�}�"6���~�m>�;D�����[)_�ã�/�V곬$�v-�9��`�H�-U�V/���_������TA]u��z�����"^Ө��Q�$�^�Y�����3f�K�M�����mz��ު�����E����b%׮�(��ґG`� �r8��#s 9�3���F��"6��qOzj��rc�=OD=lA�WyaQ�@k��2��=��%�q���0L�ja��"\���|�;��%���G�>U'�2�9�M�Z�0��z��F��zR�R��U��߃��e���/�e��g�{�8@9�02�l$�G�@�/@uc{�\�j��뽯�!��f��+'������i��q�GY#� A�\����f��u>ec"!v�6f�xWE�ـ���k޲%b���Ή��j6�A��Y}�ݖ��l]�	2��lҟ��@y一^C"�둈Yl^|�흝����Fm���u-D/����M�X@t�ңT��ǋ[���0��f:$��S%����(oB��1^EEĬ���1��[]�G_�*�?KZw�<�&1���cZ&�x�Ac�S���y�)_��U��|tC�_�q=i:�"���7�UL|`��O+c.�|RB�Q+���U����ۏh�ufGq��{
	"�&�ʎ��YY�lr&�r1��yڿ����*
F�M/20T5�<�|���H��+����jyg�G|�c�p$�g�L@g�ZLpr��a���� �OYO��V�L2��힆u-	V�mF���q�.��0oɝ@<�W�gX)ƫH���3QH�����F2&&+�?��)��UU*�b�f�«���AF�����m�on�5�X�@�U����F��.P:?,u�m��j2����8L�n�h�n� /�=��#؏�:Q��m�K��.���o��em&Q;���GW�d����\s�ْ��3VGK[�O�/C�\Yk���y��O�-:L��������E��*�8H���nS�-����:�7�ʙ�Wj!}�,���D����zP[��sq�P���lγ��ʑ������ܴx��W��8��dn�k�C��m�om� ��@"���$K]��z��S�~Uɛ�Wz~0�؃����<QJ��3���N�g\���p��ؤ���l�����X&�w���bt�HN��hD�2��4m�c�.��
��%�U޾乽���L<���v֛����N�����I�`V�5�W���l;�O�?�.�U0�%0WSE�7my�жg�qw��d�L��a�����ү�sp0Є)r�/���&�%��_c��h��6� �D(��@QM�](�6��sY��"��v�7f���i�b,��cO?Sо�Bh$�n�=z3��r�ϋ�"%���局�\P�$�C{�neM0@h�� T��D
��Ҁ�Dq�����Z�ĉ�P������8D�C��-��`�q{D��&g�DۑtEn���g�52�z�����ީ5�d�������t����5:6�����Xoܐx�kz�Wž[�b��4#�L���L�蟶W;�\qJa^S��V�?�A�Cz�1hf��If���m�;��#�@���g�h3x�����-�J����9��%?��l�g���?��a��K��DC�/�o�t�ҰCs839*�3a;��2ƿ�Y�K�����WA�_�2C�[�!����#N��C�����N�v�
�Xp�Yԭ�E��b��|�c�hU.�'���uGLW���������w������5�V���������Y�����Bt϶��o�}ɤ0#���$�Z=Cr��F:�6}��qm�Hf������댶��ˉ�-�R =ld��)pD�ݥ��h��Tp��߄"~-���`���hl0輅�)�a����eBl��V?}G�R����"a��s��f�&AL�2G��F�ձ;M��ɚ:��j�i����b&�!]I�w`�˯_�r�tݹ
���)�ϕ349%0�W7"��%��֠o<z�m]��!.�<���0�}�Ey�]	4'D_�ߡ]M"��f*���<�f�:����	Ɲ4�q,Y����E�)��������hv�5h��n�������ƿ��#M�
��)\xW�3�T��&͜��]>/�
�bBc�|�N���
v.Q����݂U�AL+j�^Q�NIln�-����c�{U2)�������+�W:��f�$���㢜�P��*����$P[���O���h�堕N?R�ᙆ�_wv(Vt3�OO{W����Wߤr�I�|�UU9�m] ��^K»��^:��˗�	<��+����!V ��|�Aí��*S��D���m?k2w��"��9�g��yόF�gQH��歚�<�*N����v��9��=�\t�gn�R�n��M@���k�+�ǟZ�wt�I��ڂ����ai>���B�x9�1�lh�q�^�!uE�{ff���C6_EׂM�G�'��������벫r �Dξ���q�8[��8>2*>�o�|Kd�my��"�`k( [f;�G�&!�T%��K*x?�O��O.jrЄmfW���DZf�w��>v���(l���
w�(!����:M�@�|�ܨR-�:@ R;9��3���h@9��+7��M�D6���;�V�%�����<R�w��Zi��Ȟ��(��s(��/T�oB�oݤ�������e�xU�f�
��,|����U�������!QBl�JV�~�� B�{�x��>�Y	CC~�vM��P��S�$��￝M�(�l�W��V^��j�G������q�ӵ�5s3T�";E3�|�i�*���7����osBIm�	�8IyIL��e`�@�9q�Χ����%�Q5�B���a�X�r7B�����)��� {ΝY�g��&�B�
m��������g[N8�U��Of�ɒ3Я��+W���8�<��;D�8�/�	}֜�N���vM���Ӻ���r1�S#��N��U����F��s��28�#PO����I5(�q�9��7C*8ԡi4�xz�&.a���
/lw�κR�Y��&!1J���VM��K8 R�e�N��b"�9i��C�u��L�F���h*D\H��Я�{�Y��=�`���·؊`����>�oOM�5K�ib����ɭ̔��;�L���00�i�0<g^/��5������Y� [��D-����eb�g�� ��7wO�a��lͰ�̮S3��k'��a����G6R��Ta�W��DQ��?�L��y�QhP.�����%1���Dz[�L�_�Qk���C�yL��a�]a*U���W�S���'�\�\�=Wr� �u�$�MC$���O�5P�]�h�)��N��r��@���K�PMC�,���?���{Tgy� �9�V�V �y�_˒�R�6R_@�1[d$V�Q[�>=]���pN��s����ޛ }N�l���U��,��B�AU�l�#��j����ߢ7ao���@�P*}(|��׏�^�mv^��X�M7T
��#�����<F)�fW0��7q���Nl��0-����O����:�A����t��7�Я�eE/R��Ļ ��DhHE�-���Д/���A/H*�5S�UJ=A�7��r�	(��CœvW� �}v�g�YPI�	+�mt���yxˆ[0.x�3��D3 ��`�����A&? ɉ�PS��4�G9�m-����e�wO$&�80�<F*�ѵ�r�YZ��M�#4����N�Ʒql��U����F������"���-���a�Mo�~M��=�f���^h[T��F�B)�+DLֽ뼾�9W�a��$�d�Z�մo�����K?KsXlxVHYEB    fa00    1200ir�E3h��$�w_g�3���=�4t�I�^�OqQ?m��d"�t,G��1`v���%2[0�5���`�g�Y���pD�H�?�6��+����� �H���@'�0҄�"Ʌ�*-9kW����Ŷ��6_ϯg00���_��>�� ��&I(*q" ӗݽ��M.��٬��f�a�v�8.�A���={SXE�!	;�l.4�,���4���"��T������/V^#8+&�F�p�"��]�E���ĞH(�#ēCL��ޯX��+5Z�� ���O�x��Y���$�`o7/0<.]�� �ASU�y���$MFʐc}>�$�P�J���ط�>�����9rI�����z43�z�3 �$�b��P�#���i�6��xzE�c��K�9��+���1�-�&��%#����������v!+����کE�t
D�A&��u\�"���&� W5"��[7�<tO���������D��R}����	u�3ԧ��d�S%*�ۄ�$y�蛋L�a{D����˕�?�mwg-SfNqƮ�#��:�Z�%ME���=��җ�`ȱ�7�{Q�?`�8.�f����ju��[,��L��,n,;����j V�����qV��_��]�BV��N�P����'�tڄ�I}�k��k�*��+.��,�,;FK��LT;�M��~�d��
z$q�a���\��;جT���ܕ�c����O�{9C��������H�xx��B2*���ܞk�zZ�_:��M�
�e9T�`qT�J.�?b�3��˄�c���^�i��q���u�º-���c�)��������ɂ�'����Q�, �܎)GE���%X�F��k58B�����G�I:k8�h4SK+ GB�<|X}.�7'�����h�m :�t�w��qz��tQ�Ag�:�q�.�r�w��	@@�b�?E9��=xh�v~v�`6�爉_��=43�g��!��0ﲡ�Z����a$~ayk����8��[���@)J�����/�Έ�s���B:	l�VEv���a6�q$F�z���IZ
W��f1B0�"j���R�ᆣ�1ӝ�.]����&��d`>߇�,y$v���naD�<��{2�u��5|0E7[O!J������Ƭ��RĎ��ƃ�sU�m����{�S^۞���=��^&Wa1ܽ��B�q�{�~K(���3?�-�;/vv�o�j@�M;ܗ�s"����h���x���ړ�W���_ .�Y��0�Twh$B"���$�6��rF�O�}J��>�璟�͡��+k'>�䚆�_@�nhQ`#�BW3P�)pXD6��UN�� ���̋Ȣ�ġ�N����eIͧv#
�p˨��@u;��u �{�T��r��Gܞ˃�_�r�r� r�G����y �Wp:`��(���/�~)�gÝ���ٷ�sֵ~E�D�'��G�GY�v���!��K��ݹ�ěoa�G#�� y���T������tmQ����%&�Г�[���?�j�k&@��؋V����޽'3�)Ef�s�w�E�x��&7w ���BD|j�׾����y�K��R6i�4Vr�u�a��BӉ�CAY����/װ���b����qsS��}i�
�'y ��#�.�Ef4\�����6���, �9��J�Lj�s������_*,:qY���$�Tf<msd�-�4�//��+��փ�^""^�͸���Ʊퟻ�!�%�qSldA��vYM.�S�סw�yZ��l
�<���`���gs�A#���B��n�����m�"z�=��ܥ�i. �X]��H�6{*�,��;/�q���Q���V���d_�E�Ͼ��e����ǯ�Lm��G0�lO#�t�&(�2Mo��hI/����Y���⧪/��Ŀ��`).�!@=��q�[�X�䎽kB]nC'L[}�X�2���ku<>p�!p>�g����7��˱�We?Rr��W�c?e(�GeIn�d�᎔�}��>�֘�w/:7���ǦSy����Fw�)2w���P�V���*��/��g��7bl-w!� ��;i�(�K�e�mE�|�<����U��yo"	뵣�M���s���fѻ�����l~rz�g�@zx=68��~'��L5�)�����g�*����Q\�Ʈ�A+Q*�7a��Ψ�Q�hj�;���W3�@�t1��S�҂�0C�������1rA�������}V@g�/K���H��v3��䡢�av�N�����}ׅ�q5���>�ȍ�g�ة��ur������Y<����Ȕ*9�Aa���Xt(��=�TD���|�~İ* @�A�]��&�=b��=l�랳Yl7�5�@�q@&�(x�����<:"�)��1��S��<�=^���2؇��$��Uy�u�&;M��k��FB��=��@v��<��=�z�&*6tJ����z��p���ph!}�nF�))��X3���K�ܨK��Q��
��[h��-eN��s�Cm�H�D}E�^��°��wg���ʵa���zvb��B4<�>��%R�\Uq5�9�,�����^
�rn�^��:�UM�[�2L� �7T�f��B�Ƀ�;1�u+@QO�S�u(SC'M���n��D�v����H-C�m|=�}��v�]�R{���v$]�s@϶�l{g2~ۚ�u���.�Q`c~��Md�ΨM�ZV��p=�j�>���YR�uJC�B7��t��}�7�+e�2ªAvh�m5�$0��U��1�sg�ϝ�kQI�+ojR?f`͈�"ln�����i6�j�Z��;�Y�bL����/y�]��J���%�NS�l��o��[j�e��9xu��剏�5q�>��R¬i��r$~� �l��������r޻.P����.L�F��p'�SLK�ʈ���l�'+P2���B\�2�%�ve�{HW(5q�4�ŏs��8C�L�L�[|U�c�����e^�7@-;�����U9b�:���;�c���K�021���7�F8���V����������g��+�9u��I|LWf�� ��`4|���yv{�Ż�U�u��E.Y|*�k���祥L�'��0�&�m��bɁp�(�yJ���hx+��Nv5�Iy�ɠnɕ1����ɳEN_�΋����u�){�b���,c� R���撛���ѣ����8�O79G4�{�5?}�x���I1�^eXQ2[y�%��-b����V|(&d���l���ѭAN/�_��}T��U�>&���lø 3�u��n���+ c�px�n���.1*���r�-��U���&x:��M���Y�$M��W^FQʕ�v�e�<[#���V�iV➁g�`3�B*h[�����6K�f3lG'�*akDƫ:�3���p���g�rN�l�e�Đ����a����_v8�ު�u�|�Y�u����P�-����c��z���oh�Y��S�ݗ�5{a�&��q�*���p$�d~�w��t�G�X����:����$�~�O��g��7�x�Ah�;�@�
��H'c�	�W���*����M��ui���2J��)�pQ��p5��Ѳ�'���hGF�����ۏNHy*�N8����,��xV�"�n}� W`���sF�����\���������*I�%��A3��{�Yp��{k	c���MN7����Jf���mH�G|\��J{钪8��>oι]�8ZZ��:�ױTI?�v��Y�nAT���@T��7������!5 af'��l����v��*�γ�;gz_�x΢D�g�f~��u2|c ���I_��\s�Z��p'<�ҵ���4��;fs1A�7��:%i�O�+N�8�WWUR#!C�mbN)�R�Cଞx`�o-���,����ě��M ��1�(rl|�A�fp+E�i��$��������F		�ESgY�E�㦷C6�?��p�4�W�>A�Զ"ߏ&[E\�̡>PNҦo�[1:�ǳN�#��;1^��K�#��ʾ.�}(������6@N.���%mm5�z�S��%��gT&�0�_K�O�� p�@�j,Mލ�V^��y4�X��8�7ې��<�f�֚�/��/��%Vб�L����<hF��1#��C
���[dV�2��<#\��:W�٣�A�p�6�A�����9�,6�%��~-�~�[!�?���E9�Ǟ�,�O3�ZR�x�K'H�:�"��Zᏽyd"??�%+���2u ;�:�sSGJ<������BkR�r�5@�/Jg����_ԝ��ǿ��:�p��N�[_��v��jI��JkT�G���'l�MV�:���U����Bp.�t��x�s�:/(���-'�K(�w��2$iaR��`���t~ՙ��*vp����ց�o��e�`4{�{�l�����e��T��I9�
��'e��n�"�7���:ZL�1Ĉ$b1��5�T���_����`���E#/ѷ�"� (�QE���4L� �4к;n�*a�������z�� �ɟ�����T�$��d͞���ҏ���XlxVHYEB    88c9     8f0�8P��� �W����!q�+�/1�\`�ݳ#ʸƈ�\Tv�8BqK&;��o�^>�KBĒ*sr08�\�1�Ɔ	C�D�D���5�K�����%r�`����VB�Ku���<�hM�C�Q��Hm��Al.�E���z��aD#0��A�U�Į�ϋw��\���Ļ0M9��F�ʫ�W:f)�4��<�{���y�X����9kP]�3h��˒bAn��pr���/0���������F�3F���L/�Ț34�&�8:g.���=8	�ze�H����b�[�;|
�K���v�}��#������ɭ�_y�j�ٴtN��3">�}��mT��Ҽ�	�2e?�P���8��Š���#17�V����9:�,�i`$�<�*�l��U����@�PK�I�W�@j(�������U�$�0;���Z%�Cl��n�A��v�4� W������8��0����7�4�)�9�-Ǭ��Xqe�-��1��=	&T����D1g������\M��gh�/yb�g���n�/TN�w����0G�������)���l�oL��w��m�o���so��HUP���gC;2X�ͼ%@�����S 2e�
O���nI�+�NN�V��qWF�S���X0��M��[�*����K���벫�@}�����#�=/S��,d7�.��d�|W������+�:�/�Q[��/�?��;)����P�@�UT�ut�(�@T�"}~7_/�Ep�-E�"�֒���"S�מ:YFQ�����K�wjFE��I��s�%;*]�p�?���h���>-=�����e��;/A����_��uL}r+�f�%���gk`���=x}�8����f^�V4�!�����(BL�>�<������_�p�W�e����0+-�_ɍQj5%���>���TB��Q���g��NVB\KsU���h�M��uf���#�(������K�^J<sT���U��ȐE�P����[-~
י5�����R�_�wCq�$ǐf�q4N{��-V����	��Ph�����0;��a����v�ƺ��xA	�2��x뒊�od��t��q#SN�>�7�<M\�#����i3JV����@,QX}e.S��I��ԲZP�vʭ��?B�y�� ;���7ʃ[��Pr9�3,M��tF6=�`�s�o�����{}&�/���f�����������Z�C(�P�qB�p�f℻���x��V:J�������p-�g=_�'�I�����1>Y_^Z���$N$}�L���"�l���D�7��]�g# *��I�vܼ�܁�U�,�ڹˮ/�)'bg�g��KZQ�r��x	(v�5�����Y"ٜ���"ma��'$�Vl��yr���N�ڣ9;H��͔���)E�jv��B�.�x�0<ô��0nqP���Ș~���7S��?�PK����P�l��d9�*���O,Zz���{S�;Z�q%�x�YO(.�lYp�$���Y&�G�
�����H?X*I�y�/������x?z�����'�Y~�D��&됭��8L��4�C'O��W.g\}o���s��xjb3hs1 �����ŧS�a�ȗly�j�(7	кo�Q��=����nm^}��\N�u�yxε�����N�a���}B��-�����P$���t��&�>��M�����.h����y����L:a��x�&�]�ޭ������9.S�^gX��=4�����+��LX�_���8)?�^�W�p~�
�՗�1��K`�
�õ��yw�.:���<���0�^D���]�^FO�lC�����"aK<b���vR٦����\0v��i,�E�o}�>�io-��~L�L�ɿ�m�-�~�.�Tq�kC��Q�Ҿe�6hT&1(�z-,��u��@� <r_��X�Jz��cc�Z6c� �AM�%}tV��N��ٙiv��� 	y����y����/��E"��D�S��+�rXp,�#����W	Y�ZtUY�T���s����AO�I�LL��iN�@ņl�����?p��e�f۬�A� t�	COfD�)3:%m�v�I8C_�������Z�g.��2��ˁ�j12�6��R���C�������v}���T9�ƺ� �R�%�v�腿��*|b,E?1�F�]#��&��������bߨj��PK�0�����j�lz�	6N���A�4����p�eI�b�/��*k
��2)�2z ,S��3��_�R