XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e�������_⤜�Z��ɘeR�����8SWdtVM}�훻�cDv��[m��^:@�y��d��]�#$?����Lr�u�K�ڻ�oR襅�ߢ�Pϭ���ڜ`�J\Mb ���E����YOo�IE�=rx�ۤ����3x��nέi�ƶ<N��UP��9j���{W:�x?�v�z���@7Ȅ�n3���?uiD��0�i�$&�T_lP)n���_��54��	���������<1�.�2)���\��/�ZC ���܀��
:�D�����N�s��H�{0��g�����n<H�u�T�I�H������v�7P������>��1���	��}
FHiƑҮb/��C'���G�����qr<������+�1����h2�4��z��H��a��i$�T"��Q3fa�������Ǔ�,��.)ͫΦ+m{�*���`-��ל��)'Ņ��m�/�1Dr�� J����E�]��oE���f����/��*^��P++^�<ԣ��Z�
&��"�UC����N���i����=)+#r�v���DHEu�_}p�O1��1+='ܐ3�~/j�\�:~���`R߆z힏͟�F}��:�*�	2�I��T����G��x0�e�gx�b�k���(��ҷ���Q�w�5��Ļ-� �QY.)Z}��� �Რ�������5(J�0��C��
�=�:l��ՑrYP~r֣Č�B�ma�)q�t���K�z�A1XlxVHYEB    1802     830���/�V�S�^�ֻ?��%���E�J�O�m�Ȍ>���*��<���#K*:��H3�"��DP:���������B�L{�l3��}��h��J��ec�ƈ����~�@�W��-�!i���ڋ�_�GW�� �"S;la���#�^��u6g�x����N�8���o@q�M�\6�]��͉�ݏ��C'
�j>�D��FM�'}�T�a�@��˟�U���2���!nL(� ��d@�b���znT�4��᪜�]���s�:� ğ%&�P�.�/���C�IY kM��������?`O����%��ud�	�Fz��?D5P(e������Mp�Wl��,��yfWWт;W���X~{���D�T~�V!	�Dִ���쁀���MC�+�?��f^)8-��2b���-��5Y|%�|:B~q��D��D�TV'�aI��T�E����f���y��0�C� ��� ��&��*�D)-�t�A)���E��_�4��[��J�k���/ܼ�J��c�e�%�g/�T�_�l<Ƈ�}6��B��"��>$>�ø^�n��V���]y&IX��Q�j�xu]�G'ht�����w{���4��pqr��BY�u��V��r��,:�[��Dm�P������g���?�鼂-DA|��NUeu����^�t���[蓃��/RдS���'��:#|�)71Zy�{��MT�ۢdB�}AЖ�g�ԥRJ���K�7���� �7�p �"uI� �ќ瑶�/��%�;Kr+��lA���rw�/t��gq�6ס��BTϥ'�Z��z���ѓA%)��N���Lɪ:��J�)g���'����f�����[>�I����OO�J�ء�� ����Ȁ<n�jk��D���o�0a�ۺu�uX!+�ؘq�rpU�b��饹�Y�
���@��C��MAl�/�J�9&\4�����!Hн@����<�>e��s�$�Q��R�J���^#�xMup8��e&3�j#e��7|g�.������Ϭ�T���8�|3J7���w,6kR��u9>��	Min�|��U܄�7�v|�_K-��A�7�i,R'׭�@~S}��o���
h����C
x���p�Fr��v_QCc������&^��R���8��c=���~�s�M8a'<q<�H�}���(��ω;�?i��"b��t�����F<G[�1���2
�Q�n�t':"Ad�eq�7J�_K��͒2b�����+�0�pD^ֲ�"�?Aj~B ����L �B'�e�ϊ+�BG���e%,�F��C������]T˵w�D�GSV`z����.m`�����ˇ4�.ex5�%F��b���_�a&z�F�ubK������4D.԰��뛤�I9a�K*o��;#��d�
�$�h���E|k.�X��cd�[�z������%�������`F
��F-��$?$~���)x�3��n:�z0e���<T;Z�#���:�5{�������4�Pd��xE�/��{�����vc*Η���fX��郶8q�@�ͮ�(�,tD$��@c����N�7��w���7�]Bk��a�>�Ƶ�FZ�"��4���}�V����l��	�E�a�l�!5
Ϧ?ڻ���1E#Q����,�����+��I�,�+�Ӛ|n����ԕ"�y�}OG����)*؀Wo�bmF��oO����b���)��{���.���ǖ����9�|}(�4��W�Ԕ0��0C�?R].���Jô!���EB.���HCw���#���v�R���G:�itz!f_GgύR�k1]2�4ȑbO��j8yE��Sl����!��
`�k:�S�
��*Fr����T2s��3��x�'ʇ]?������fȅ	��Q.�7��Z~jV]o�2a�����?E���7 5�ڙ��)i�@a��)�����,=��"ex�3�V�/F�K�Ǯ'S��z���,uc�q���`�/d��O�	�6�E7����v��ʔq�+Vvń�l9�Y2����
z'��?�J�_c9w�