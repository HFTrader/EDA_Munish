XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��bW��'��k���Tbe���P����jv"�xyW�,{h�I�[�[�.��ɍ[�oeM�2���M��L�t�t�5��#�D���g�!(��UA~g��`����>&��Q_��?e���Y�|^��w0%aO�j��.��1�`Ȍ��W3�q#������4�&���&I�q�+QJZlp`�ق8�y$R1��� ����1�v�lXz���#_���vvI�4P?�N6:���A����hIv�8�B���<�0� %G�oil?�q�?ګ2���Sq�e@L~v,n��Z��Iy��$Դ21��bW�����I�'�Ũ�6����M#�{�K�xR���aT�;	����<>]`[��
o��
-�J�੻X�L,"�XC�s$�KF�(�gh�3Ls���`��#����I��4��0A���pdƴA���}#��u��١͹=(=���	�;�O	 CC��./��#K0�f�O�'Ud�a��R��!���cE�4P��>7G{�nO0�s��zw J��;��o��-�|$��F+��7��D��YK�����F4"�0i�K��i�2����^Z�D�v��Y��s�|x�5kH��0��вx�̤���բ�����A�ݣ_���[>R���h��o�ŽB݇�#��+[�� �ԙ�϶h��B5�麴�u�YAܻǒ�y������`�-�����N#.�_cú����փm���5b��.��\�cF8�/�ًT��因/q���2XlxVHYEB    160d     7d0�J�q��.
%0��ai���9�@#K�,��O��η��m;�=yV5.?��)Z��0�H���GC�"E�F���!ڋ��%#L�NsXK�N4~^�!;��G�YWM��.��¿�u~����k[�Xf܅�~Àc���ZÀ��iAR:Y�d	��p�C`�)i�j2]���n\	6mS�c���4��~(����J�/	�����Y��Me$-#Ӌgb���Y����hf-�]B<=�s- 7b�mcAb�Is̑��8:+�ZzC1[wHF��[�J��c5�۸.%/����Z�:%�����o7������qk���b��}rp[h��&��֕��ng�>���e�Y�wZ���ޢy�P!�_����o�8�!�"9NC\�B��cꈺ-�>(��ݺ0<�k ���;?o�Z4\J9�@C�!�&�):Ȍ�[z���m��4j��{�0�%L�	�v2V��P/�Ru���G	��g5�`s#�|���3Gum��������dcM�ϝ9�u��xz�{[�
�l�z���g��M���Rv�x���U�Y���2^YX,p�3���!���U�9�,BH	�`�k���
��b��uh��Β�){l�u)�qE�����*�e��+���m-;��A�#Om�An�!6�2!�^�Z�����I��f2��8�O�$@���q'so���<=�� �bBf�#�"�G剘������G�еnO��N�NY͸��/���q=ym>)!yl�oQ�N	U�4I�C���M5�#e�	q��sS%^�J����}X� ':f�X%l��d��_�����3���(�ݸX����m��K��w�O�s����I��o���\�2��rHn>8i�"����\D�)��y'ct����m١'�w���h�x�WTy����k$ P��ҬKc��H�� `�Y]���&���|J�Pc�!X�=O�5%4԰B���vE/��C_�~�&xȚ��?A�/�X'�N�є���dY\��H?#�/����#�N��w�a/���(�+�̷`�
ԭ�E��
����#��DǏ|X�u荨F��ո�!-F)�r�����l���!Rw�4u�1ȈB��I�4I�#.i��ozNu���f�� �T�k~�혂�F]�w.�"[K�m�ƣ�^И�xQ*��\p7z�̍���S��O���Yh�x����o�l���Qǰc�3�/�_:�Gi���mO�_��M������7V|��Y�������sࡿ��[�E��H�x�\˘Y3��~��%8��d�?3��ߎ�I�QS]�6�fN�7~�ޱ�Ő����ø �X��g�{4~� ������ꩰ!���Ln
J�+�S��5�7�:Ʌf���t!�`��m��  �NfnMC���:ל�>���g����lfpq/���.0@�(ڪ057g�لu��j<ri�5�O���p{6,y��N ��K��E�V^�h?�?���5��S�c��	*��w����;��;���[�A*n���5sߘ�U�yw?]����;ސL��+6�+�g0-zgnQI��1��8��I��n~�rX	^W[9�N���M7p_�+�����������Gh�G�q��@���д�+)�W���Q�ܤW�{�E�I;�*7���Q�s4#��7N�D��U������S��Q�ui���CŸ %S�՜^�s��^	���x絞PX�)���QWabu�a����뿇�l������h{Ny6�9 ^a�X ����K�L?�hG��GY/�$q%�zD�As˸�(�t��B�|B~�Y4t<�������0J�N a��.��fg.���w�ȑB7��H�	L!7������H+մ�P.P_:��8gs,��aْ�̵�x\�%'��J�Y,�;�+�#=T
�z��(3X�`<�Έ�^��[Fn4@�����$^Za
��j��p�f��Xu�2i�����߳