XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z/.��ҒE;e��q��&I���\��!��@)8D6{��q
U�´�d�0npDH*�����1�KBg 	�Qp��6�b���&��{p�9g�^�V�^p����� �o��:�VKp��7�� ��f��eG��!�V�&�Jp��9k�0��\����TͭcJS�@�N�I���ָc�Fh���AF�����㒾˰N]uCM�q�����L!����%��1Yp��"9Q��̺��ɍ��L�tu�4�­ ���a�������o1R��o.p�0�'a��o�}���.L�t���Vή��gR�A���Q21�NQ��@c��S�^�u#pǄ�~�i⥲�9�+�̯����3eø3�&3�V��_ �1^!Qu��Fj�R(%�Ӏ����Şw~����֊�<)��i��;��C�v�����T���X[,^W��ot4M�d��a� yE�UjC���i�~�.E33�m5�yEYn}�?=3�0A}�x`����]8#<ύrY�`:���tIţR�9vi����n"��]7���e�X�v������Dp��gA��!)17�l>?�Bl�����lY�s�|�am��p��E���{���/M��v��)�y^Ή�|��}-����l�%T|�L���z���R�48��٘�ׄ�R@Ii���Ix";+m0pMoӯG.Z�=�������h�ymz�UT�����qk���q��I�Lv�h�@��6	����z;��JG	1XlxVHYEB    b631    1a00�g��Q-��VƇ����1�pv�����>����|��i���ڰ�,oj�����_<d�`�3��N�[��%T��,��5GU��B��V��mnZt�����3x�,fq��	�,�t� ��T^�N��װ,t�U�C������h7��R3�r� ���@�HҔE����bp}�� (s��h�Z�{�B&�\@�l;g:1.�G�%���^�&���6.?]+N�p�<���R�
�@1�=�NݴP�c]�� >�6�ts�y�K�]l��R�����}i���!�b�t��P�,��[�0F��/�o��MX�M�i[8��l�4\"�3;���э�c�-��ɒ>Ky�+~/8�]s�����#R��8���$e����Js&Lv]��$[O��1��4]� ��Fn�5{�\�%���j����n��������$8I{��(�����"� �>�*�liG��S���/�pM�Э|B?�����*.�v��jiZ&�4=N���»�v���%'�Z��ݿ���_�L_���4s��zyo	
t���\�L,����<��9�w��g�e�T���f5�ZȉS_��ʫ�Y�yOR�y����N�VL�Ce�S;�N%���������4@����v'�������/��m�M�i(�"���u�,f)B�����%I?�����V�z�8�<������Uc/JG�r�ڪ�W��3��H�q��L�/`�>�b�M��%�:jH����	��z���ce�A����W��ra	h��Ø5<j�S�-�O�ݗ]Vt0o�9�l�<;�Us�v2����d�����lᤲ}eʈGuV������`Ɲ�2��%�A@ �F���	lw>�[�e���26D��~xp&�Z����Z�/<�y��P���+�*�y��������E��0�>��|Y�+i-M
���!��e�-UӢ�56�����7�-��}Ur$h�!��6%
���7��x!�R�~3�!�u�d���{��WN�J��d�L=�4���(�:.��"�`LwR>@:�(�N�s���S�o�5S��n�����e���Y�ȚA�$>B��ِ?�N=����֙,}p��ȎdO}�S�_�Ph��D�(��ά�P��[�����v���7V�H�hr�{t��槐��E�︔���>��՜l\�Y�f�HN��9�J�.7v
!MV�IvZ=׮�tQ�� ��f�Avǝ�4h��IL9c4�f�b��tg0$�)"��N�B�F0��m�p�7�2�碒b;3U����9xS��'
���W�(���_�/Ri#�qܜ1��;�/{W�u#w4[~M����叧�wa�Q���(�t#�S�[b��U��:D��Sl�bD�
.�oe�q�sL�f9_���2Qn�oI��9����]I=Tv­A���]Z\`@����T����Z��r�6#���{j<#]��w�ꭞN%,�>j+Bc��+���~f*`����^x�V��|HL��W��߯����dN� U�n$�����(�����M�(��\ʘw�\|-��;����g����ފ��ݲi�ĭ�t�4E� �+B��������JB����f�NFl����0�:A��'^iK����L�EY}�'�%
<'����%�
�/3��1��;)PM+q'P
G��+��l�!a�l�I� Ɵ��a<�XR��K���LC�Y"D��@��ƚ�Z�f=vV��'7t p�^��G	��?G�*Sv����]�3 Hc�,�?h>#7[=�c��6�"�\V-�{	Ǎ�܊�}�^]�=��f��)�t3�c��Ƿ�.)���тb-����t*�AIkQ6Ǣ�k)��,rU��&G������\�g��Tz&�����I�:}$��^oƒ���}���4ˉ�̜�����-qY�q���"���UwAk��v�>�i���O�j[p#9�+��9ZPA� �ǰ$�mi��^[sݴ��W��̣\E��/p��ù��>yՎ~0��V7s���2�yp��>��©��ӛy�9R�,�;y ��[�E�_��	?\�YH,���ibh>H�%�nDXF���j�K���)r�DT�)�^�غ����F�9�C���PS������(!?:��
};�$(ږcx�8�pIpW��]����"�D��:M��}�=۱�;�*m#_���t�W�B�+k�~�wQ)�0?8��qj�wW$:/�QҚ�"@m������3{���F�]`[0�EG��'��)��#�}�<�`��FͲ/Z'��9jE)<&%nl�ފ-Wv�ӊDy�m���cOnV Պ�Ȭ�a�
4���<��eaxo)��&���+��'��_�p� ��`�����r*!z�7�OleK�Hc���1�lm4>.n;['<ỗ��0�"�������dw#���=q��I�"�ks@qmb��F����?� ��������xK�����o�>�dmZ&�sg�<꒚�z<�H��j�7D� ��]�,�CC�y��h#'�������a�N^��Ni�=�װ�i>��f������C@>	��-~�<\|�na�a�:�G�;�9 �5>��&"&���,$�fD��fOxm�hR�~�b/�Y�dl�&�"G�\�y���WmZu�A��j�]|ل9D�U��L)B��-�/)�>
=rBE%g������WU�a]F�j�1��e�^z�`�p����O���!O���|;�}��o�Gy���G�!V5e�����O�� Ai��k�Z�%�����JB���#��@-��5�6�e����|�7�+�-�K�"Z -�����7�+��c�	a)���1ӫs����yf�s�Qq��f�����5}�zQ�kHx���G�L�d� �n��فw�X�0�z�"NeT�ď[V���H������E�Cn���R�rڶd�&fM;?9c���[̂��!�$
�����vQ��������P�bh�}����n~:�-mz�����!Ӣ�� ��B@�"��)�D�����1W�ŹJ��	�Jک��+�*�5�#��(
Ȧ�G:�d���\|��� 	�x�m��l���|FR��&�-,ɥ�T��\�"{�e��a��!X���%�����o����V`�Ed�Ҵ�ʯӉ�v�%!H$]-N�-��4���E��KVǳ8bEQ��_�/�$!o��_��
��-���V��|��n��ިRlH]Fs���v�g�@%���V���~;,n�{J��RQ��M�i�������LwI��|��r�����l
�HR��0�|��Bޏj&#Q%01�@�Pаk'�yP�
%[�sg�{�c�A�(�3t�r7QE�Nc��zX�*�<�$��d�2[��Z���/�N1?Y�1��E��@�9�>Z˳N�G���'�g)7���|����#�j��Cv8&&�i�uZF����,(��(0��e�uڅu7�g�<��"���`����:���v�=���S��c��!��Y�{NE�[��p�8����ܨ�;F�ĺ0Y���̾"PJ;�zpqX7�%-�
\7��d�$k	ׅBW�״Z�0�|^���R;�#+Ay�H��	b�@��������g�h��+t_�sR�g���\*v�&iw�'e!p!)c��@N���FF��M'-��O�:�a�u� >��v&xdsM��t?^��`$9c��Ջܖ��FY ��_�ڽ��-�s,#ҧ���L�x�+W���;~N�Ei���� ��(�FM�/�-�ޮ0��}u���"�F��y��3=%���T�Z�O�<m߼��'�:��)��כ�Cb*p��B�z����q(@���N/�JK��F���`�k�FŷO�.����.n�DV�9��s�B.�\�����C㾭�ݙ��|�@.�mOi�Ӆ��ۙ)O(�ϐ;�j8�f�X�\�&��M�_��z��
���I���j�"�R麮�ʯ�����}�1@�9�U��v6+�ЌuY��ԡ�X�;4�� ��Z}\ [l�f<٭�R���q�ͺ �O�:US�������(���4�sh  ]�oU�ng��!�T����� 9N��W�>>u�zF��ܯ�f��}�֖ ��}K��	^	�S
���{:�Ι
;��1�NAQ�1/��Ff#6L�J%®wf� �.%��"�~=n����2H���w��A�h���oj��/��d~��0���
F����}rD*��U.�v���fw�F����<����8nro��=�.uh�����+B �)�}k���ro��
(�sʣg�@mnf�̪ǈv�`X� ��}T��pl�[��s�i�"^�3�OdH!EL��1�:��_4r�A������%�Y���DX�!��2k`�o4��s.2]�
�aL��$R2�M,Cᢟܔ؟��n��	��ś�9���L=<{o�˄������]�	�d�<b>�̒���P[&� ���S�t�j��>>�5���6ۦ䋒�ϯ�ʀ��F���`���!9B�+F��N냧a�O�6x�+"�*s\!��>����׭.%�|׸���VI�?��4��@��,��'��s r���4ϭ����7�P����2����7��pw����T|U`�Ug�	E����F�0OڎUT;z��6�  �6���k���ކp�c�:�]�� j�������c��A��5�=�DF���~v���sh:W(aV��S�rI�_��)�@�
^?���h��J�u����ht})@����(��W�o�z�ݗ=�Mz�٘�8����l�	�bit��;{�X�$�1ۻ�
���r��l�ǎ*n]7��MYש=:c~UN��_�xB�elzBz̛���J W5��{�ğ�)�mGR"��e����.������0�K:�I�c=a:�����'ti�@%UU��[�j���z�0c�M��:&�rk����pX��x�b/{���y�l����� �צId_�;5~ii�ª}��2F�{��}z(մXk�ѫ}6�(�����=#tt#��$h�n9�,#���ִ��D��)� '�{�`TF��w��G)�-�}�>�0J���4��z��D^���cƔsؓ���BW�DC�'T�CK��sB?Ō*����[vbe>�\=�';�r��t����UM�C �1�Pd��O/&Į$؅��J��|f$.�
����A^�)F����(E<r�ݦl�@��( v��O����'�>��4�ƈ�[����A��-\�ۥ���%*�y@�Rؕ���3�O����)8��QF�H��{h��1�&�ϑFM'R���7�.���3c�%���?�A�Λ��D����S�Af�� �D��?ܫB'��;"���C��h<��:C�.�<�D���З4��+�I}4�����.c���2ѧ1��F����h�P)�M�j_��K���x��x���-{�L����g˲���5�Lʣ�'��Jx�7\�(�$�橩7�H0�KܦY5S���I~>��.�>�Sq˧����0l�#¿=aԠ9
Mp��u�{"��\�)�c���ݖ�ܹ�9�3nJUc"�Z�0+��b����;.+�I[��x�aEV�|�u]���V�>�J��L��gSʉ�C��H�)έy��ʨ�V�^�b�'O"E�GՈ��OZA�!�7�'�+:�U�������.N�;�ԥ*�^2�(���Yɩ�\c�ә|�{ł�������X�ڡ_7b6�=ڇ�R;���#8A8��Y��߉���{{����Y��ئ5k�GRv>����"�������OGQ���t��C���݇��9{+EF��v��:�)��L�ǅ��*��7h��c������te���a?�b!��g��د���A��)���>da��w�Ǔ��o��+��(�(N�{�U9Y)�iV���6�T�(�*q2~e[�ӧ�*�PI�i��o7QL����灆X�7�u��.|Ᏸ�o���Y-��;ZI�-e���Iŧ�1,}}@d%��$�e������w ��#�_�;Zla��cF���g���S�͖%��zϒ�֑̔�����S7)�;��
1���fK�� _�<諞q��+��z� �i��Z�L��"zq��#�u|fl� ����a
 Me ���j��xe��#ܱ��<�����C;���g��NG_���V*N�D4���p����"qə|��N~�S.�SNe�����`�k��X2���I�GZ���K�LXo���OW�꿺���T�ȡ��J��O�^D� 8��b�x�c<��F��kr%�}݇��}i�&�jAb��T6ќ�.]�Ă���1E�ٻ��w: �.����gR�C<I��K��^75[tQ��m�[�͝Ɋ�\�]`z��Xk(��Z�~����^��;hg++�#�,p$����g~��-uYS����l��ȵ�%%�=LnJ��$j}�܄�0���:�q�J�0^�yW����3�t���=pN	=�؈qs�t�'z3q���ױ���W�D�8�$Z(����!�M;�\