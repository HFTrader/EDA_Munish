XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���uz)�#��A}�~c$�r7 �<�'h��Յ�p���D��_h���Q�&M��vMr��|���Vi�K��~�A�*tiB�"�|��������}���\�o�Փ�a������v��?��TW*\E^k�A�ᙸh��Ȁ���|��l*�֝�Rq���u���n����/9� ;���S�6��Oʌ�t�G�#��zܽ���X[kd��"/�'f�t��M���&,
��|H�E�T7���)��Ou���du{QS'k%nU(޾b�GEӅ=P�K,��^,�I�h��{�����:3%��0ē3��Mt���U�@�G[�g�d���G9O�ޙ:`���9�o�6V�՟-���Ƀ;j[����T�u?�a�<͡IG��2~/G2�S`����dzZ�~�
[F�[6ո�Gœ^�
6���бU �\��vD��^|ΰ��=�{o����[i��WC)�J�i9��*'t��؆���`V�pm��n���7A�ҀQѿ�p�o���W<gUH`ǏD���PwWɱU��^	��4�c�������E$Vr�h�І!�>�N�����m��X����S��vRrL�ﱑ��!g��"c?nK�G�\�K��������g���4�M.�����o�E��t(�g�� �Gqh���fӰ�^�X`��^m~���CmÖ:dS�m��fn��,Uip"��<ϩ�\אն���&�'ʦ�}���f�[9��[EN�_iu�l%{]�Hc1{0,s��XlxVHYEB    c6d9    25d0�OoS%m���I��4ٜ8�&%W�Y ��a�:�'%M�Ӿ)�զ~ìL�6�U��E[�<�!m
��|>��+���+��dgח%V�[|� �7������)�~A�=oͭr��޶��@��e������nd�[c���_I�MMa/J5����3����xk���.G������Ą�\����-�pAp.9�o<�Z��/h&���DW����P��~�Sc����}*te`xʄ�������1��)'���lR�s���x�p��9���3�� �C�F?TQ�]E�ZW�[PϿ��Z㯐.�wgjR�\�͔`H'��t�;i'���7�5-� >Vk6���5�uc��/
�����M�*$8NTT����C���ys��[oD1�r�Ol*��2o�8�j�#^����A�6���/C�j$�#��@˴���dh[S�D�2��������/8���$�8B+��Lf�$��fFD\�(L�	���i�O�����B=ه�N?ɔ%�Y�]�C*]�h���NA��
y�ʞ���[�/:]�]��Ʒ�r��%t�<0�b1�n��C��{衲L����pC�\s�v�x��r`Kv��M�~]������8Nb�'{I������v|ѕ�/��a���ѮQ�
@��'���P|-��n�F���/�����f��oA	-�~���R9E�q�e�Z�Nv��� ����6z*����aE�����H��)@�O����d�D�����ݤ]�tr�ϭ/9�㦧�@E�����,2���aejU�"�����_�/�1(6q���$��ƣ����'15s𥵄���&�5\���l�:�C2��)�c�� 8����ӂf�[�4t���S</�O��߆!���2.��n�D���d�t���Rr5oR�!���Eh�+M�������2ܿ���H8�,�k�>rb��? % ��HP(����k��z��}ki�xu�N�ʻ�JF�~Y,�Rr�$�F�Q���I��6��U��7�|�c���t-��?QE� Ŏ�-A���l*����p�w@"�t���.^��(�V�����ck���4~��l�7)�&����#��9*�t=�_�v����bcB�r
-ia��V`Ɵ���Q��@�����ۻ�����NT�Jp
�tԧ�W�U�Z����Vh�|��������~	�����f�5��@^����U_��at
�~�,W��&NR�0�[���-�H�*\��LW��=D01�|L~t��rZ�a�C���{�f�~����;�TN$腉M���:�E��t	|� ":4ݼ��W�5p�xpO&
�l�S�����t��r�T��rݛ��JC%a+�U��bp�6A{�Nw��s�8C�5�&�.g}��£��HǏ@���f�&����x�:x�q����QH��.]����ɛ���~\W�$�7`�ĺ9���������K��
G�y������������X[Mrr���ƃ����l]�χ�n�U'|h�:%�<�Ӱ�ӻ�J���k�h��s��މ��h���d(pw�J!:gm/_��$?uo�쌠IW˴��T%�)�-7 �&.�U̜��5�����*J���*���ʆ����4?���¸���U�7�����&
=�B��۴^xХ?E�U�L�,u��ެ����o��?�g>��D���
~vLq�7|2��Abi�g+1�D���O�3�)7��O�3u2��?�W91�F��瑧z��UV3����[k�7r��M�֔��dZU����[h�����X��<q�X�?�On���R_��*�zp�O�D˵�`ma��Y����[O*LU�̆�7��)tv;� R
��^�ֹ����?e���j{P�7$���'%?��x���i��Ӏ��X��R�_�	����T��0������Rd7��10��՚�>�>~DK�MJK"�)z�N���i��3D�����n��"#{�o���+�|R�k���f"��[�2�%�N30��/��S�T�SlB��S������OG�l���|L�"��}�� ?	k���L^ʹOQDj�s�ܢg=�BqXm�Q�>���oN���RǷOK��]գ�d��ߴ�M{��vAo���5�o7OG��'Q,No*Xu����2���./^�ۊ�U��o�zA܈M�nnj���Q��@쉚��m^���i�;�T�~ �V���];����w���H���8?r��[#�W
�mFz��[��)_��}QQ𭊖pY��'LM����b��|�H�'ײ~(�b{��F؄�_�T
���x������n�18��_lN����^k J�$���C��|��=JB�dJ�f�j��>������դ���[aUֿ�-aP�������;/^B6�}�����Հ-ܧ�[��ѽ}��rS:v�	�a������%�z�{����@������P����a���ƕni�(!�Dκ��0m���>^��)����~ӫ;�H��Ŗ˛�giU� ������y�mXښ^*��w��m�5��il+!4̐]K�����x��s��S�(�U���������I����`Nu*9݊�h�	��-OzO���\�y��s������V�c�-����m���Ve�t"D�&_�v�:��J�Fs�L��l�iO��RV%^�Od�bn�Y�!K�|��KD*7��u���x3:a�RlT 4��0��� �Y�j<��ܺU��h�D��qi�9���KO�t����I�'O]�e��<��dt�zg=.\ T��䍎+6mI�h,.�Dq���+��1!nԃ�6S��B��k��&㮱شa�5T)������56��D��_�c���l�zu�V�Lz�?���kN��R��8��1���F�g�6'I��1�v�w�4bi0� /
2���r�F95cGr1°�0^���Y-��=���V�CW�w�IŲ�w�֧s�jq�@��B�C
W�:'Y.�R�!��}��[]�᝘!\8�����j�\��lw���:`N�-k�Cd��h���D\[?c��V �Z�L��)��6ΐpO��kB��
-���Ѱ��A���E����֏�eV�nj��~p��#kJ��U}<��Z�ʉ��c߻Ɖ�l\��	n�W�8��BړG�m��NQ�X�3�m#���.�P��P��xl<�yO�YG�I��_F��S���充��g�C}f�/��۳C�j��~[z�D� ΋��.X�#IB��WT.Z�)ft1;��*�D�Z�ȟ�2L�km�~���s;��S< ;�$"f����m���e�-u!�riL�k�$}��~��?UL�l�76,�1{�J��{�&�T�փ������g�I�>��C8�h�������C�m��� ��ik¤z{W��Ʌ�f�~��cE�_ʣL�7.�Ӿ�ޣJ�	k&(V�N�hSX�2��Q�����u6�?��*s�I�&e�a���]�,H��5F7� ���U����qM�����L�����R>�7��x�N[���Ĉ� eׂҼ��s}�wU�fಝ�l��PW�I�'ڞi���%�䮹BЏ���V2��N��	��;c���	E����9��xN�Ab���	�c��k�F[`���vV#1J��Ƿ�!( j�d	��U�m&�)k
���aJ�����t��.tN*9d�"��5jwx���L��4�&�Q� D�
/�k'���)�:��kuv��2Z¡-N-�{D�r��Tlgnr ��Gz�{����엸e�a����ҋ~��9#��JH+���A�G.�e 5�p�$!����Q�����T�0�04+�)r��eJ�y��'�18`�?�&J.9e��?ѽE��hS�+	�G���9�4N|��a7}=,�ɵ�VF�ոx��>�<���Rey�OU^��W*��\я�ȵ�F���!	^C��/�(�|9��f ���X씂�P�&��F���	
1�����B}y���J������zT�I���K���	���N��E��J��*������j	��⭒�@� 6fn���,Y�K���ZuJތD��Qs/�ƗB��=�ޮnqey+��h���o�����x����N��i�0��~��zţ	�-@F��*��^��L�5����ݨc�,q�M��>�06>�<s�,�:���g飦a,����~R�����jZ�S0�<�`��v!�����w��Y�+�t�'�|)����`5�H�2�(:��?�(8�1oW��0a-��_
q�.���a]7��eT˛x��)�f�L(���H�sh/`V��~�� ؐ��.�0�q��_������_<~�u.���`$L�@n�:[��z?��ܲq���,�'	?3���%3�c`��7�ID�N���{�j_�&��}��z)ksC���6sS��mr���NـC8j���rZ" �0�F�L �5!;���袶�qb�}��i�t�o�t�L�����`E�詼�+J���th�9���������=��ޣu�dȭu�]%*?�=iǙ�7�'�֫n/��_�kpagɷfܵʴPܼ�5gr���JJ+"d��>���7v(vH�<uf����A��K�Q��!gK�]_�<\q�7�n�!��� ��N��q~���0Ԋqp�ӖO&�!^��fO̼���c���|T����lx�Sj��!}�fجY�)2kOZ�X���Ѿ�k�bhu�e�X�v�_�����v'̄���ٻ��8���{(/u��Ƽ!W�������tB|*�����ގ��cn$� e/5���;�w\o����X��z�i��iw�$�����OWe:��r�U�Ѫ֛��t@�%�?C��u�'<�l �@U|�>b��*jҥs]J})<��T/bH�vw7�_�}'���ͥHf���o��j�r6�7�rh����v���tۓ��9/dy����G��}�|�X,H|�ߺ��3ҩJ̘ 	��]�� ��/���w'�{׶O���J$4���8|��y�zke��Q������6�mӲ�Ƞ�}�׶��51�г5�Όb��-Dj*�6��~�M$b�r�:�g�8h�Q�w�
�,:Uck�<s+酳�V�W֢!���J�\%�*�}#����jW��rş��J�y��8����/Վ|J3�{Rѯ̊���'���I��ʱ0(�.�2��))��	�s��u߿%�%�BT��%o~���ݕ��f,ӽg�]>Lx���}��糦ሓD��)���(k-(�rXt#�'}J�G�iG���~2R/{Ť ��q�о�AqؑۍS��l��"-Tnxw�����;S��3��׽A��d�k��)P�1�X�1By��w���	O�b�b�O��אcT��� ��S2G����ғY5���%AW�*-
�<�z��]On]l�c��1��vC�a�� �}��i��y2h�3!�H�fʊ_���I�Z�	Ay��sS/OE~mm�f
���DdD:���sX����9-�"sM�c�M�)C�!e}	aT$�+���J���L
�0O��ū�`�iI���Xʤ��T����
Ԁw ő��Ǘ(�eE>�pl���t�~�G\:�=>��M��3���d��7x&'�<Q
�&О�y��v��yѥB-������|�$S���+�Û'��T�B^���=_K��-�<W&h.��ߛ�t�^~)f<5<-�=��cUV�W�����R���~���8�1���¶���y+��'��n�\;�c���?�-��|���V�l	A���cb1�e����бH �P��e���(-��pJp� ��L$��jF|� Y;?���ϒ��3w�\>��a���II;��$Td�;�}��	��q,C�W��*@3x��qȥ���h���a_��'��xy~q��`���D��M�zm��q�9�.�U�V9Y���	����2�|������+�/�t\=��/���_O#m��2ٿ���"����7_w�l?�\��\�=��8SQR6�����6���U�)�խ�hp/��T����j�a� !�&�.�PN5�Y������g��j�dZQ~���9O��ٓ7� ���
`Tt �08�6p�h�o��x�X���B��R��(/hH;��`Q��)lD�)b�xO�ݠq��Q��P��J!���BmȍJ!N,�YZ��v0l'Ke����1�G�y!m>�Qj�%�����_�B+7�q]i[�,�;:r�³�]Qy�~�h'0Z��>@�f��/�J#� �����`ܭj�p���
L5�vL��ك���z��r�[��+��@�$>��vF�;�����x�?G�7=��X"�3������mCG��Kkˋ����~F���B	��yv
tG�v� ���]7&����0o��ZiLJrg-h�*D?�����)�_{xi�c�H7w��,�f3�)���	�S[�*�`�+PF�)V|VJ賰TZ%��e��4�0-,�#���Z��z�J�#�6���I`q�0�7-/J7r�e4���=�N�v��rGn�bKe6�x�)4mQ
W��b����n�\݁�y��̑a%�m,�]	�������B|�l�ܷ�QU�'	n;�pYk�,��[�T�V�j��|���ؘ�� �%�GZ���pˠ'�X���EyQZ��t��#�:�W:�����+�[v���P@�N_�<���b����}��$l	�)�����J���KooEX�1e+��4�E'�(JX ���ޕ��a�j6��j��ymR�A7��k~�-'�~u&&1Hց
��j���и���l��8�9󛾹� mW㾃�(�7_ fڞR��͐ܖQ��
$��XZ��:^�_����ǭ�zК��z����r���WE�9N�G��?�hCǲn�G��0����S���;	�y�%�|�8@�PS~�������� ��,v�BTx��0-˜ZJ�C�H�뢄�7"X��m�a9�֬5�\�)S��A�;�7Ek�lH]?���r�8@��}w�w�8-c/#N��^��y�:��z�����
��vw4��%b���xӯ�{�[�Vt�t�t��	��D �De����a!ba�����t��q��l��gr���Z��u�"��6� ���$d&cM�>��|B��;��\�9eӴINK'C+�����B��\4hX����{/n��6B�kpxň�߆��l	5�Xq���lp{K=5Rh����PH��`���;(]kF˿ub��RQ&z�ל��y��_
)��&�A�l��ex ݟ%fg�☊�G���I�:������`�5sq��C���c#Y�*Y���$U��!_���H%_���჈j����|��^��S�c���pEB/�.Y�)+n�� �VhR�w<��b��h���lgc�R���7�r�Nl�`]��1�a���3���.졟���[B�Ias@au9-@�>�űw	P3|X�����%�*}xw�z�H;di�V~�����|�7�B�O�V����ݏ���d,>�1�<�/ڻt��f�ѐe�2����]��k�`�Cc	��h0�-8a�m�Q����hj<T�B���I!�3�$@����Q�8N0oݯf�ל���S"�,�8��oݽ�=��S�&X��%6:��J����-i�#���t��Ƈ��t�)�5�ۮ�2ĺ�z��]ґ�gkc�f�B2ڒm:ሲXf~�'Ϧ��V�������H��g/�_͓z�Jj�&D�짢�)n
�(�'n
fo�ָǮ+1L�!�������Ho��J�k���7��W�U}�7��b������lW*h��-�=l����vD|e���G6s��M�����������0z\�D���0���<r�?��6�s�k��
h{Ǫ�h�����ai��C�&�Vv�=���.�*��[ݍ*�[��xEF�	������#>�˔'���	�����=Fy��<i�Ȏ��D����p3Ґ����[��)k��F���O�­˻��)���)P��DN���%o}}�t������W}�,�����`�֋C�]�Tq��m�;5�@�E�W*�zZ[ /��[|c�4�;�q���
n3���OZ��6��(�b=t�~H*I�Ow/N�p���=��J��d�t�@���Zi0�,k��?e�1��;���b�6k|Iz)�}�ԛk�,��;�R`8�wL����lx�^�b�fد�u� �).�@F�U��{�K3�fƫ��/��&J���E+i�_ ��z�w�8��mUf��޹~s"��j�I���<=�]۠�K�W����Iop+��
8���2�~~�t�$Qvx�a��%*�d��v�:�>���r@ˬ٪FHP�!�N�\�D�N;�Hl�Jw���!i�{�v����o���h�?�1��<��W;y2�8Ib
�?O�/v�GR����+��ݜX|���pkl�U�Uh��b�:��`h��p*��e�t�sS�ը�� �vq17��|Gف/�R`W"��ն���]PC?]u�/&����hp���f���(��c�1j�b�71���dF,A�����2P��N��v.y�"���}f�H"/LR�E�=7� ۯ���� �Y"����(l��`x�]3fZ�����sC%[e%�[�F���-,
S�N5�Vü�Q�T ���
^RO����7���Nۙ3�3I�̡��橣
 �ܟ�9@i��$�}g��*k��%�H�$l��AA�#���k��ʜ�'p��D{��!_w�aoe=��1f�r{��M�PB�<ֿ�\�����0�*��VNZ� ���0�@C�g��r��і��՝��O
I�)݊ǟ��Mh_��#G��T��R�����#r\�~Gej���A�V�CW6��Aoc��DCrzs&g8l�3���v18�O���'F�U��oGX�6��A2q����+7�TL��b����H��}��V�6�F�p54ت�������`P��7h/��O
J-��i#�ގ������tgy��
��9�k��sb��d�k	�5m��l<[p^�ʖ�U���z�"J�A��|T'2�][{.�]Z��02�8�p6���'@9o ̤iN�J'�	mՉ���'po�e#S$�A��a�1�2ւ�Z�_{b�����{7Y����半A%�rT>��?U,.<�2{N���K�F��AҡA��[��bd&
�����EkV RG�y�;�����14w�������V�U�Z�N���Ⱥ��=�3���Vp���+!��d@=>��;v�|)3��Kd��5�Q�p��\x�*��%ə/	�鋇l�CN�l	����k��e����m̋�ia��CĄM�(�\Nq:²��B�{mH	�N^�������7��wA)ג��ߔ��"Ћ#�����Z���@�Fm�\��<��b"�/�2F|�����R=�5B�6>1{ĩ+� �kԖ��EO(�X#v+��F���!�!����J��`R����#��s��Q��\`��b3��zJe����