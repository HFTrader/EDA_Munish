XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��f� ��c��%����V)�h��W�sL����lV�`x�c՛d�=�N�R�˃ϡ�ieA�a�6�������A�P���:�����^�D���l57��7�o���|Z�GF��n2�ˇ�ϟ�P����0���q@>��6�KvBopZcScSJ�&gk�9��%�^�'/�8�N�}A���5����ʔ���z|j@��g�Y�DQR��9k�f�P�^!����%Ɣ�V�S�=�D:^��]�ƙ�^�(�B�Ϫ|U\����G��K���C�"R�u֫�+#��FDM�[N8f�Q[e�'&�p.^X��:^�l3�	$�'~�G�'������V5��mN�����Z�OT�ܺ�h�C��$��R��.]*�F���%���@[�th�&x"��JA�iv9(5�Ã���A�0�4�d�E3���;�&���xQ��R[�|r��S�ƺ:�+3�$�~(~��F�W���e᎜}Պ��� o 34���r��j�H�fF�O�d�l�4�� ~#��דP;�]@_�_�;Z�������I�_�*u\w1�h��H]v46>�N�&�ՓYn��g��BT�S s5�yco�"$����,�>F��w���lԤ%�>�6�{ �R���8����Z~BlAX֛�8������C��!΀0�)�ۺ�F:��	=�ߌ���ܯ�/�7�A\?��?T�(:�bƷ����p|A�)�����HI�Q��՟��0qu�%1����@�6+�����XlxVHYEB    fa00    1f70�),IJ�c�[��J稃�箨�-�;%���)�����Kύ����]^�g~�f��p�ɡ��8:��n@!5�/|�q�~s"�+��%��n��]_c�:3��qf�7�0mt҄�eTƌP�R���0`M6z_��rE�r�G�2Bq�:�轴Y��P>�_�\�cu�̎q 3��O��dԘB�Ϲ�]��[`6	����R�}\�kl�x���g؛�IC�=v-������Y��P#�7"�2M ���0�%w���[�e]E7�4^�U}��������wՑ���cմ`q]�����<�[Z;Aخ`Tn�]oE��^WW~�����S�(����4тJnh�L;z���sbd��y��+J�%��:�}� �$�+���i~r�k�f�7(�$�-��W2�ԌbiV���l�P�-��P+���xV��,B31��]U���b�O�&��y�@�&��J���⡶��[0<<��������|	�/�м�l�'9	�|W��Y$gyӄ��A8��.�T�Z���YG��F|=��q�]B��?0�C���f�#�A�[�>���i.��t�yP�攆��p쑟w��O�A!��ߗ�����{t�S���u�X�"Gq�װ��8�"r�v��K���Y4?Γރa�zě#��Y��D�i*r�D����IƴK�`P&����WC߸x�+ޗ�6"�G&"�	� e��v�m����tH���0+:�#���+ꅪ�7,UW�]�p�\5����'�R�G����Lx��Eg��Vk�>2;e]Tԙ���:��<^��Њ�鏈J(]����6�М���V�N��-�b{0�>#�V˲#k���3�ϖ@)d�ld�KA��,KNɬH���I��tL��,��9Y�N��gD`��fQ��5���"Gx&��sE3XŘc�Ju΁H��j,Rb���L5t�9�\��#R���4r�65��c⁕;��A����1�����7	R.��?�~�x�<�A� M(K:V�Gof�D	{D��'�'�j�9�E�f�{A��<�Yd'Vf��^�p�Oʔ���9�w�6�m^{Y�V��͗����񮙉�8�)9��CZ�ZGE������D�D�rpB�:Ų�{}o�� "��_P+�����/N�ׅ��������f2�D����H���.}��Gۄ�:���"C.��%ϲō$����	�Oga]�w*�xQ�����Z|��z���xN�6V~+>NF����,2��e�K�2񱒤B���gA!w&ӓ�\�j�R߫���[Q�y��@��M��B$^Jes���$�N��h: 0O%��t�)!;N��AT5v���Aֹ#�@��Q�ڤ�~��L떋@胿J�ɖSھ�O����/i��,x�`�*"�k�&Tr�Ui�7>�ۨ�⁁���R5���׺΢n�Y�:�E���y���ՠpw�<X{8]1����мӜVP��� �o꼕�T�b׈�<���M�e���ZxD,��\1�;����a�G�IYgb�Yc� / ��S��@Ͻ���t�s>Et��:�d�1�=�C,SDIo*��q�v���GM�}
J^BI��0�*9{�J�'dn��%<�=�/~�%c�3J�o���D\6��~;����LO()z#��Z�el"+)��wV�% <V���t�%�gڦ�ZN�輡S�-���5��28�q��T�[$H�J3��,��a>Z�e�Lo��{T�5d:��C{;."��&&"z�=f���j΃L�oV8f��:D'�AS
&�R� ͎�Q_�<��/~R�:@~��D��$�ȓ��̪f��j=�XNe)�Sr��LOX�+�6"6g�g��HGЪ��i�w3ܯ�=�6��g��l3_�g��s')y,��+��X�lP���ښ=��U�Z`W�������j��P��ךXr{�GU){Ι�I�Gl�2ja+̬Kd PX,L��գ�t�B�4�s�fN~v��~o�Q^J�(�5s~��H�e��$�f���������v�4+vK���#�'�֥�5�]}��U�r���i�}��S�1<621��˳��P%�`�'vp����KC��aބ�x�Z��<oe@�{�*�4�h�"y�NxQ/�P8A�yhc��}�����/'6�r��?�����)�����PG�&��p"�-�nt4��7�E�� �w��)��)'�kP�^O�1l�;=�9���邂p�F�Rr��z�m	�}N�k���<!�P��������y�3�8�2����A��6Y�/Y\�s���6�oj���o*�M���w
�z��`���4�e��o�����)%Aji.��X܌=h�f��o�F��W^L^՛���Gh4��
��=/�a1k�vY�"�i�do2�W�N1}Ve��] k�gj�f�[	ec�8�'kI
�-�i�1&ؐ��9�}[_����j=��F�Dp���WsX]���ާG5;�UVW���� �ǘ>I��v����}J(��_�?��1B�@
u��vWw�+�_�锏[�gAT���ӱ�q�_v���+�q@-N&Z���AA��3҈Gt��4�P�b�XT�S�.TK�8͘�/b�rp�.�8#8�D�=[=%�,O�2�����L[�4�O��i�-�� e����g�E|�5�|�N����q�����d��s��Q�e��+Ն/?2ElO$��1��**��la4 ���p�⬗�(��v;W�x��E��p��)���;!�HlGĲl�퇑�8eG�q%qX��}E� �	YM�i�>��d@|u��+PnT����^�/ )$B�$2z���@�׉�9���6����
R�-`Lj���6"��	�\��H &�F�{IP U�P�k�xX�/�$�̘qVL����3�TS{� 8��QP�3���K���qªR������P����CW���V;p�N���F�Z�"�vs��ؕ�tR����w/�0�,�5����Յ��gma� $z�twlp��ѥݡ�F���t��~�U�����BO<����ҭЛc���%�[n�2��d��SS�>�>�ò�M����������>z�Uv������L0t쌼^ͯՃ���1܄�H���~��T�p�~��y��_v邳ݻ�#�ʘ�C�݂>@Z�iީ�yV�E�3�[L23XMm��p�X�:���}���#�k��EΈ�H����n��q�
Q���m?~��BZP=�&ai����ɏ�$���Mn\p��U4[͒�	��/�}���/U�a��j/ӶI��|剏�eќ!�˟��=3�[fewMu��8��af��n���TS�U�G�^c��i{i����;9�p.7�u�W7�E��u��(�U��p��s�y}J����($yAY�oc�h#l��g�@�<�K6}'�	@� �̈́���xO ^�6�M|y�;xi�<��h΅P;o��~i��(q\�o,*�q|���q�M���.dSW���X]2�vAW@��"�z7y��"��z�ݍ�mF�:�B���1�y��d�kL��ʼ��B
�%�G8�"��u��M7��Μ�����]`�N߶L�?��נ"�UX uq��P�6M��м�	;�� aumL�X����w���Ng���e����H�aY�v�|)��64;�s�9s_�n�`���� �O���&���ҽc6K	�E���_�2����?	H�@B�Tu�0�3��<��g�����}*�kʌ��90�R�L�&X	<8����Mv�0�
��^%��|׹���u&Ԁ��-"�$�vl�[�*�+9�J'E��9��O�՚�ʟfFs�í��h��O2(Ȗ��A��U'{����dȿ�{qV
P��5�u,�u������}�؉#��E�V�ӕ�
�Ȗ����E�DN����S?�F��[�t�ׄ(07-�+ hʿi^�z�B��8:R.��1���0�T�R.Ęe�{o���JB믃r�Q�����?f�/�����**E2����c������D8�P_I"�+B���l�Y)90b0��oq�1/l�4��a��s/w�u��h2)�%��֥�S����h��Y�}�By<u	ܺ$ڒ�����i���b�)9-É�	�C��K�H�ro�O	�s��h�.Yrz[�%�Y��_̸2�v\���$�٬��Nyl��h��F��T!(q��V�0�n�s�1;wn�� 2�H��dZ�pk��Q���;K!���*1F�Uy2V�V���|�F}���&��18褛���Gҽ�k����
�9�IO���<1�\�(���38@���-���̫�]V��Oi�8��GiF��ե��/�Q�T-��jr���]é�&!;F���	�(ps��1ZⲙE�4��<�
ӊLv��!�e�i*շ��ɾ�F��w��<�O�|M?禨(�57��Ȁ�Ŕ���Ij�*�:�("��h*��E�F�T�˵)����Tr��J�v<$R�]��1�qS*Գ��2���7��ԸRs��#��C5$�G&�r^�0����d��\��~N:�Ҿ�^����Ũ�{ ����%�򺔇�j���N��4���ubR���}�ai�８�ELR�G |5R�.Ų��9PVk�#�WF��dn?�F�BJZ �ԙ�"~���73�4�5u⤈ ˯ޢCO��&/\�pAǦb%GTl^v�Oe�Y'@�͗v�MP��j����|��eIC ��� �B��׼?萯��S6���Zؗ���ܪ�e�o��f[}�-͕LZ�ڹ������b�9�T`j��D��¿�<b���{�Q��17�{��+�$��\��α#wҽ	��nQj:���������}�,��� !��s�g;v(�;|��*w�ذ25~i}�H孪� ��^!_d�x&R�Na~�V7rYtb�&$w1=ә��iE1�l�G��������"��Ό�����N9�7<���f1���s���ER/��ɥkW>�O˳
?�H�m��<�y�K&�q�x�өE�f�{���MO�H
�n��������t�5�,�{[�0t��qƼ�͞wB�P�s��D`�x�}>]Y;���*x�(h�qk/V�F]'&Q �d�x�*������~�hH���a��tU��V���3Ʋ~#���.;}���jv�g�f�߈Z��	�[9�'9e����}Y[��9��': �(@VX� �$4c��J�M��̌x��#r��F�\j^����4
�"�]`]��; �0_����Z!k���,C�@!�H��s��@��"��F��?��%�o�Ţш��A,a��[��yB����`V�K�Q�^</o���-8u�9�Zju��VpE��L@�FpF����ǟ^�H(\��B�Ͽ�J�#%0��[�QCN�K]�����L�nW�<�hob7�3�N�^T��K�����(G��߽ �(�?��G�T�t��7���+=��������fl����7���{�ԁ��T7a����ri3��NԎ,\c��~��A��<�M�'�B�Z���셵�HAi$��y(�q=�巐$��'�͒l��x�Z�X����y��2 MF��x�
|i��&*fӫW����'��/��� H��3��|o�q�DgR1��ր�����k��mJw��b#��c�p���F��{/�Ǉr����A�`�}┕��������m.��t�������}�ut,0-pY*V�ƱVq���kd{k^XD�?�nխ2���vV��;���E?�Ϝ�e����I5̥���?�;�G�%�&|1A�(W7����lEηUi��D��R�=��;4N {AjN"[��,[���@%R={kM�V(����}�\^��O��"vgGHStJ��|0-�0L"��} `��]1��v2!l�ȵ8"ę���J�/U��4]og�E�K�`�{gѪAف�Ù`Jk	9�h���]��55xj��s�͒U�׺Q�8��!��m�������-'Ny枧h2� [���6��eYB�$��a�d��7�x#ت�ZY��ΐ���h������3���`�4�lp5AK�4���9�a�@�����
1��w���)��>�R����QQ�b���ݠ�r�`��L�B'��&��g�[��>^-ٶ���RɊZ����ܝ��Ebb8��0�2~/��P�ma�ea}�����E��C�c�`!���K�vmg��<��I��gwF�pEn5*4A!��'2e/�o��X�A��t[ ��ȍS�^M�`��<��gC<?z�.�	 rKlL�t�O�\���cRcj᫜c,V���lA���*�|1?���d�;ժg���m�r�,��\�����1�t�B��F~��'�];�]'�+��	�*>^���<��g�嚯k���7�mD3/�0|�)�b�0���J!�se��o�g�I�|)e5Wև�	�\�
Â��X��p�Ep��@u�ӯ`a�
A3,r����'�Zn�B5|՗�ǖ�zx�ٖ���D�o��w��6�M��1���(�{��4)�׸��7�Q��սwO!I��u��~��-2��>q�1}J���\/IW�:L�Oc��*�3��9�J'kv�Ct�� Ђ���{�W�x�=�oGRs	 �^�곷�!�d���r�j�Zy	-cI����p(�r�h\�;�@�npS<C�K6�J�H-�$�@j!(�������j]sS�3K�۞^?'RמD6�8��J�$n�k?7��m�ܹZ��'��eQ)��W����L"��.�Ll��m��!2&�QBm���F@�X���f@��U�u��YUq�h�#����hx�Y)�HXnɕ�Yk� $}
hEq15E�Ġ!%�꼉�GpBΝ��r�F�Cҷ@��k�ؠ%HPHR��N/��A����}&U������{t8x��T��~Rj@�������t�+xR ����*~:���ױ�K�6·�Unu��0�F���d1��&���:Q��� w�������pe����ΐ'..��l�b��'�� ��Mv.�p���
ʪ:���	���/����+qg]�<�g����hgn������w}\���rf��D�Z �Ks ��y��x��[������H�=�k2�|숡�l�M�v�Yc��?�����!���9<g"��}ce����ﯬ�ҽ��f����jĺ��������|�"�ȐQ\��9��a���1�$e
S��<F9�\��Y����Om��jwc>���Yn�j\����4���*��y�<Mn9��ce	$�R`��6$e�2�Z�	�	dXt�R,C����N�1&�F�c��ɒ�d��0B���(�	��x*���[P�<W!�z�?���S�d�{�+��K�aK���țn��|�Q(]��E����#�[ϯx:�4�K�h3��3}#��S��b�gB  ��s�'JF� ��K��S��x�_Q�Kc���)�X|ɏ���@m�L���C(�ha��k9�R��C��� G0�۩�p�>|���.�I��To�|[,AT0$�G�.�M*/Ԓz�b���[��O��QQ'�M�*J��v��<n��;i�s����#�$�� ]�K��E,�&�e�\A����'?N@��Ch�v��X�"�_*���X�3H�T�����BR|�D�����J�^��FC��:p���j/C5υ����OXﾥOm41�
~?��~�bj���MՋ���nQ��JUf7^�����FҦ�k7�ڥ�Od���j+�~�*��)����U�ɢG���)��(�Fu<���w���$�{e,��Y��mT��`D�����h��(�+�(E���1d��0�F��0�G�y�����`��XlxVHYEB    fa00    10c00vx�窒��qN�W���J�y`���]��-E�����^��=�NҦCn$2�}��|!���@X�$��R�1�����w��;��ԃ#��i�k�d\r�}�$7"�v-;I�%)������n�����%����cEI�4EdzЉ�鈚�y�yD���ڻ��3��,��y���($F��[�d�G�.�!D���;c_�3F��t}~��$�G��~��w��A��<�TZ�4!/�����lЛx:3�X����q�e[�8̍�:��"\�����Fci�N��8��/LN�o��rO�Y�{#1��"f���_V�::�.~����K�s8��\M�C��4�Cu��RM��D@Y4�~]/gЅTJ�89�x�7��γ�2�>*� Ӝ� p�z��n�;��ih��Z|@�+"`E<"4�hf�x�F[җН6���W�͸!���^s(=Ռ��L�_ �6��U��ȩ���m �t�l����=0�ڣ�[w4�����g
 �D
=�8 ����z�[)�AT�\����g��Y�����>,7�B��'|5�+ b�v]U?)��pM��c�L��j�=�%��O�R��3C|TK����/7�f��e3�BW�i���,�W�:��Y���@��TȜ�VM�=�]�m���,�"�?�9�Yi�����6P�"KR��"�;g�O�����2����ۺT>���$߈���Y���߈�ȫ�W3m"	3�h��>�Aq5�{\F�S�z ��
\|���<��B�7�\nJ'�	���]����U���'<ŷ�f~�!����8,b�ĝ/g��i�\~�CF�bxP��ϲ�^r��$o*`������'-�K����>�n�*�HI��9��k�"�:P�:;C{r0f��%��N�O�"�@=1@�H���+p�<� +kl�Fbk	#\�pw|0$�L�(e�r z����)>P.x j���N|�񑵺jy���PM��T ��P i�]�[^>gx�{�đ�K�����lы���_�E�N�l���H�w�}7�.6�Q%&����75L��Lj���"���e%w]�ƫ&|�$���8������0'�7���T�����G� >$���i��]ц�c(Ǧ$�[��o��O�q�\�iuY�,U�O��B�.�$=��֎s����/Lt�k�O���GW�~)����A/��^�L�[�-d���L�@9���Q(�.;^�Ѓ~v1&���
=��k�ou-���G1zmE	/we8`��� ـ����	�����]��5��OJ��B] �����/�h��`�]�5�
N���
��N���^+�~x���5_�G���&�z�"dD���b��m�rB�1��Aa��k]E����[C�Ζ�w�k#�tΧ��#Ñ�Z��l;�6�^�V�\�i,K~����BI���L��T׍Uc�h��%���b�.T�nF̮�:��¹i�m-�M����b�	�$0���p˯�o�P1r1-�<�a��+������ݬ�6G�X2�}������o��|T�s)�73����%cz}y�=E�j�f=F?��z�-Ǧ3GJh��{5k�|ѓInVW���^Vw���P����l��:�1gB˨N���-������6χK�s��-��ᇡ�J� �� ]2E�zXz��s�X4�\�7�󩗦TJ"-�9�C�rC޽�QaD9b�R��j8@�d(�|�E�:����0���F;�{���6�Y��5!��:��ӓ��5��?�Y�6�މr]�Mur�3��0i���֑̣R�F�g�;�M��ʆ�pO~���!��n��+�K��]�]���d�(�V�>߂��˙"��� &!}!�I���Z��r�r�]��)^1WRՖ�2�b	��'����/"���oR�A2Hj�oN��=E8g��;���w��Ｏb"Ɨ��{C��(�n��n�^IلE�/�c�B+�Nu��*�i�Ģ<�ocՍ�LC�TOw	{8�W�Á�*�W�z��?,�V&���.{Ԯ��߂|�]ue����(4��_�(�$�m�܉L�(��Mk_�~�S٩n)�Gs�5OS%�dj��,���Ⱦj$�Nwt�\�̻A�����H�x�*�V*�~�D(���4�ԷH�7�3�a:[�Q}�۩�ʠ��1���W�v�� w:*�������8I�i����>@�B�]�j��hk�n�9�a�8RL�K�e��A�i5�~ُ��.UW��O�fSUqg㐆t�S�,".C8�+�zvɵR��-������\˫��^t"�t'bԐ.0��![�r{�<\g; ��LZ�����l���$��C)���|��F�����!�zs�ڱXl��v)B���<�1[Ls��k��R.�r+ac��Lg�(3�@i���n^Q�:H"1���{�O�*���P�`�?>r�Q���K�(#�|W�.��r���n��G�.�nX?؈S�a��I�6�1dϦH6�3n�z<&q>>�w΃_����oc����1w��P=���\����L=��qg��q �F��pBm������_>���>T�_��*�5Tv ȃ��*�O��a����c%�_j%�OC����*u�5��)�v�"RW7�T
����ï2�.�T�#;H�C]���f��Ȭ�&����(�%�å#��+Sɫ�N�� +Mh���������db6��+�;sRj��_F����h���4Z���n/�|��+�h�W���1u�9���MR��[[�+fo��RPv�X�+¬���3m��F%���O��K���T����v��<��Y\���ı�g�*yM��`:8[�%)N�7�����b ��f�C�*1:�C�"jr}��f}G�R��rN�����V����i<�S���#$�� !�Y�v#m��Y�c+\	M=�r��~���(�����hh�����>�2-?R��3yG]َ���M��C��XQ@�������<r�K����)hPp��X3J���f�H�A!�@�4��VY�Kgo����@��([Wy&	fh�毸���V$�d_AY5����QB_�r����v��t�w#$\�}��Ψ�t��Ճ�R�3�T-���udJ7�ݗU��v`ا�롙A�p���
�} >���r��Η�Qt���'`�<��wo=5
���<��=FS�J4�R����d�J�]C��~�"!ZR�0��O�1�&1�D��a�i�s�u��/[�@l(^��;(8���E�	
����]�_{���#���^�̘,��8��+��(ǜ�Y�>����Ә�<���(��P�فȩ�6t�l�r�L�a���I=��7��S�����7?&��9w/�P�aEG�B�+f1f�갴�f�Z��D,"��y�`�g�%��A�4 �U�d�niՎ�c��(�%Z��H�_55�Uφ��%,9��\dcǩ/0F������&mzf�'�I{�+I���ͅ�%��AKִd�r
ܗ�ϐBE��D�%�KQ�1�.gh����K�u��������<��m��N���[�O�=���nw!������)���5C�Q�?�Kp8 H�����*}�:�������Jߌz\2�t��F�w��3��Cd42���^��[愾��2 �틀:��0��׀��^��Nf6(͡S�������z��2�5��\�!O`���'�ڣ�ķ Y3������{Ӡ��[�d=`�X���$��D[B�s���^|��� #���a��k~3}3k�Ul���)�+/F�h;��GB%�DoT��Dc��a�b~��@|xo&ݥ�?
�����5�lt�C��cjH vb	�7�l�|���$��-m1|��l�����yES|��� KS��Al$!�0F�4��c�TF�ّ{Bb�^�1��@��_�*_�g!�'�����Ti�n�8X�\S�6RU������{��cg��tUh��U���(��0q�}YZp֧��ɚ�����i�h~$�g[/�x�lʜ#kH�|S$�?��b�Yh�Wj�9�pg�(��YL��)�������R?�J���~I�Cr��JM�k}�#XX��`��mt�� &ڳ�C�[�8��:ђ8"�_(��"ц�ᴅ,:l�c�o)Z�QU�hW���Q���&��`/-U�����r��/*b���.���$��2k^�S�3zy��SimLB��=�&�m�XlxVHYEB    fa00    1140���2>I�D��t�l"��bx����2�
�Y�9ott���!g >d`)=P����s|]i_� �NQ�9�6��\���a̻ٽGe��_*�l`��W�}:ΐ�b�l?%kc�}~.w�F�U]�z����e����.�zo�*���+bu��"���u�=	
ɜk�+nK>ю�#������Am2؅Y��*�i[;��:�j�ǲM�O�3��G��=��$��SF�4��-I�����2��Z��J��P���é�Y����eM=d�G���(SM��<��[P��;:�F����t>��p�Ղ�`��'���ʥ���A�rP���p�s@E?��Y}�,�J@��c�ע��[�o�ꃟ�����	*dF���Z���L���ׁѾ��>@�X&o�v	W�I��!?��^�[���Os�͟������[�R�Z�1V�l�_'j+-�����N*&��#r���$�g�'0��h����M�Ɯ�!��_fTQ&^{R��)��t�#��F��z��Y��`���M�*�y���	vu0!�l�51�)Z�!RV��f[����i�������Rv`�w�����3xc����'!�S�7�P�����%=�3��}=[�r���y�2��K[d�
�@����Wސ"����f�~;�c��q�������U|P��Ɏ:l�.�R݉u�'[.:b���P��c���T�(<���ּ3Ma#I��N�x:?����yݣ5-L�X)C���OcN�ݮ�*�	��t�?͐L$�l}o��p#�n���X
rQ�
aX����T���Z���xxb��K=,lmԻ���I�F<4ק�Ϥ�	|xF�<�٭w���e��0ھ��5�]����H���m�6����cƂB��zZ:_7N�ujy9o��1�̮�w�4����Z3��1C���]�L�'�h�s9��yɕׂ�G���=��b?�W��w�&6'*�T�p�>du!I.��`�R�� :��G����E+��8�Ig�2ɒ �F��n�	ʤjT@�C��B!}\7*��)�����l�T\��_�~
MC 3ʬ(��|l�4���c�8�nǚ7/}Krʥ�z%1�j]�E
��[��+N�G�+�V-��]��=�Cr���)���닆��N�W�"#c��I�2�%��*�퐫:3����'��O\,���R%��4��aH銬�:������0�=�)�q\�2�n���M|��Kb8���|���0i��Ǎ:����~��#BK\��/B<�e���������Y^���E&�"q�+;0?5w���s���uex�6�.���c�93>%P�7�χ�jt�M�i�o�H"pDC�rH��ބ:�c�ˊ���Lv8��o�T�%F�]�])+��55�/p�Y�TS?'��2����	ɩY3Ǻ�v�U�G2�H�<<ZP>��1*�_m���b�P۔�Ўq�e�m����f���f����ˏ6�!�A�#z��X�IU�p_)�F ��hC'q�T(c \�÷���d>�p�̝-3}E�Bh($���FP%ѝ'���5�����.������8�i����2�9G�
JD<�||���vH��pWa�;�G�z�����6|�h�T�|F-!�~3�m9@7tN)�[�u,+�n�����iC>�����h�$B��6�aAݒ٫���97\WK���u�;�����j��s)1��4������8T|�o�˔��;`fR"Ý����q*�Sb�3�����R�V7�d��Y(�$��K�hn�C1 x����Ѯ�E�B,�֔KWkE�0�ŵ�0׈euJQ��m�7�՝�Y�hO(�ZB<��W��T$'3S��r��U���H٥�i�#��c�q�	�lR���4s��)�,�S�b�LF��Wr<J9� �2�z������MU���t��E��H0��2�W������J&���'Z�{��H�P�����n�QN@6݋>�GQ���hz�g>�!J��Z��v��f��5��k礝�uD� ��;[�����x�'G
��n�il_AfJ��X�[~l#�ֆ��v}g&�>�Rkϼ�낥RV�r�fd�Ӻ%�R]ꅵ�ϳ�F�ލ-rý�Z�K�0���\o�"
�bɽ�3�PPoE}Xl}+���R| S���
����kVVqr��0}!E�X��55G���7�o>���E���/���G�����z�o?����{m���,~>��E�e%�s`�n� �\��oƏ��g�E��sr&yQ�m#��E���4��{_*�n��/,���{��jE��K��W�me����U@�O5d�^U��0cX1L4��[3�Sj+'>Q��R�CRsp��k5����ϯ�~8$�4�Y	��>����9��g�4��\�O��Wr<XM������$sn1�������/��z;�M�hl����>U�_��F�"�(������h��O�Y�;�
b�	ZLs�����<@�!���
A�R-~̥���R��B�LZ�cVi���>O5թM�[��=��]/���l����2�Q��}%������%���[aQUZ�h�F�$֬��i)��U)�w�I�F�%�
�S۔�-@�_r�}z^��#UU;
d���rl37]	ci
��#�rID���UB����sW1��D�c��������ȃS���[$W�*�w��7w���0Q�'I�(��>��o�CS��^l�&�Ğ�O�#94@�$H����k���`�Z�\a����ы`�_��V�_����F/0q��xWq�7�^j3�,��K�ug�.=>�&��ɸ83ۀr�!��$���q<���7�]��]�>�x��ng'H?R�7�k+�jE���@>�u�w�B'_�YoA"�~��Nߪn5i��3��4��:���"m����H��a��ߓ�ڧ�6R1}п+��^SJL�k�7�)c����IG� ����S�BD)	�U$��A���K�ZBB��p�ؚ9��k����[���{�?���.>#��=��z���θ������X��Z�J:�n����F&\949N��I���	�fҔ�te��D��
f�� ��=�H2��?�u�mft'^���:�>���wl/&Rx��]�M�T�;����ı��19���V��C7�i�:\:�J0�Y�]#'�7[:!?I���v���~&�3mP����)^�-臞��.B�_���r�oInz�����l5l �_�o_�޹K�ZD��0�6�mz��J����5wظ.�D�c.L�oC� �\�W�r���pf�kDT��B6���Q ���4͊�'�J*Z�{Y*��`T�t�}}�f���4�g�4��,GK��s«q��Q۬��u��H�f�`��n�O�6�֞��(��[8"F�2� ��J�H���ё��L��g�\�#:���+�U{(�pD5�j��шݷ:.���Ldulo��HǒRN�o�a=�"�?-y}�Mz���D�L�U��)D9\Ӳ`R

tm��t[�x���D���G6R֬��47�9)H���R�@�,�1��3���z�W,�Z���\�T+g���c�*k7㶛��?H�4#0�s�� �2F:�%��u� ����K9�P@��H�?��+�ܔtp1������lɫ�i7p�!P�D�臯��H�ȗe�=����z4�O�.�Bx�F��paߨE�䘣���R���)¶���i>��� ����CNHtpCpU���8p�����@�t�$A�^6"M
<��I VcF�8��`���,� �� �)^�5 7���¡x�/ �S�`a�#��!_��F��}AUŖ��[l\8p'�>f�\����L�rq�A�zC�?�&�iT'�HBb��9T��Ϙ���u�u��[i����q�:[w��1��X��^G�*j��F?4�[D"����hW('OT�޲�^Р�Վ�Y�q�n�>�����Y�E��MP�2�S��rPo��1"��B�g KmH �i;䬄�\�z|g��
��-�k�z֥)ԊV@������|M�H��}���dl�^%��ٟa!�q��y�c_z��Ѿ�r:јWr'd�dNy�X�|�v�qT�_�C���P�`���An2�q�غ���#3B��y?ʔf��#ZCƍ�2'6�����~tӘ�I�}꾩�Q��l���}�)n�3�1c,l�p�5S©��t7ESi��k�9!�5�� ��[:�YYk����r��]&E�i����4�Ӧ��:QJ���N�Z�m�ߐa����~�9zb��=���qg�o"��Y~�������Z��5�n>�g�D�bXlxVHYEB    fa00    12e0�+�c��V�O�T�%�Ff�ߞ۞����7� ��Y4��	�$�K2i���H&��'*�n�*/ٱ�[Y��ߩљ�6�؂i0R�I� TyE�~�?-��Z�Vg=fX%o0%ϐ|����"��s�����q�3j�H�$ֲO���(o��-p�~m6��e�+��]s�ܼ���-����h#red����i=0�#!S{,��K��C��[�b�	�%K�`C7���F����g#�T��D�� 3���BzY��+�[�ܽ���صX���m*ɛ����2��m�觴�=|���
*8v5� �F��	Gu!`����t0�����D��0��/@�.�m���M��d���4�����/�,�Y�b��U��Rî�Jr�s:$0O$x�k6i�9�m(	S��$@ ?�ŋR��9_w�L�v��/c��O����3���1�ѕN���9��v�̶�n���Y\���;���6b��sk0����Q�$5����YL��J�,�s5K�dڑ�C�V2}-].[&�Ѓ')�vDR��ب�I����'�)�9�7) )0l�9egr[t����B� �&�*l�����%ʳ��^dh����Z�ٟ}ېA��T�[�N�_0�`������Y��Q-�ȟ��=aC����eoQ�u�-����b��c�Yt�O�:�u��B1=c��5��҉H�7Y�"��C  �h����u��R~ ��\3iU�\���3��eČ�e���1"͐�t瓄`�?3���!�@ҷ�l�G=�(�� ���ٹ~:��6��6H� �&�A�cAr�����c�c��"��T��"�D����qM:���o��T;H��q(0<e��Q���̼L�_���o�)O���������Њ92>�]�� �L� 8��"�	�����~�X
��;�Akg�x�n��6�8ňl�>>3(-���b�m��>�A����/��7р�o_�>��*����t[���.���]��_y�s�r�vX\w���ڤQe�C>%�ܧ��8��6z�E��4�M#+H'%2..�4�	��wT��bշ-ޣ*��khR�L�cBH~M<u�:���W��'�\�d3Dt��	�~�5���|9D^Ö�9#���C��}�B��(�6��x�U�G����D���F��zԽQ�.����o6%� ��{���ղ�7�@��]��+�~D"[�Y[=I��?�����+!�V�w�{��T�/�~��C(_�E��ߖU�\����.&4-9�
�?_�;N��8ɵw���	�סz�1(��1N��´�fO�������Ә�m/i�|�f�5�����|ר��1�E�_s���qI�6qb��4�;�`*m��5MةQ8,!��� 5�3��p,]_ңO���̲�{����Ѣu]W�=�:b4��X��t��oYƱf�m-ֽ�o�]t_(|�}��T9�4�9�r�y�ȳ���-���3�b8b6��+���M�hX�AO�U	��BOL��vY��v̯�;Ӊ�8\��Q���H
�~<uI+xuU�0 .fO��i4�DM_������v�^�^�|�o�����p�Z\�H\�Ϯm��ߊ-�̢q��+).�QW5>c 4������}��V^��mT4)������q�7�#|pY	˚S�u1���P�]���q�䖍��8��aG)|�X�yAz�rJ��4lJz6���s�s4�1�t�n���l��T��6c%G�F$�ޱ����p��B�e���]�ç��3��!�<��cq�!'^�|�CI,(�I��Y��K�Y�BA���mɝ=�ԉ�ز ��`�#��k�"�cྥx]2ң��2	t�qfy�@�4��N{���I��Dw|�%��Lڃ�}EQ���!@@[�k��Ec��Aq���C+y���q�.x$�ap��J���+� )������\F�Zv��H]s��I��ӋWOp��\��k�A�H�v���'���1A��h@0`=?L�N�2����f?�NBD�uks&Z�܋;b���kΉ+7�؁f3Z�RWqi��5LƚA&	����f�Lc����o���A��1�ƅ he%ơ�.�L ��p!~�2OS���V$3 �����x�(��J��lR�YB��޿�a� �>C� �W��q̅�;yq�������;�}#�4dG��ތ���C��-V���5Y�,@[�T�nf�I.�OAm�!X	X$��wa��7�0	��;W�;v�P߮̩��+�6sC���d�0�C�]w��h�����$΃̔ˡ&�zo�T��M.�ca�_����#��I�x�m%�-�Ri�h�"��nے����
�/0�j��|~lX�E�	����O~�Z}W�q�T��KP�|�����h(��+��h�U��54}k��8�֓ ,���J�~c�e��EcPE��'��(�If."xh�R��LJ\���a��[���bf�v���Ѫ5b�8�Y�2�N�ӿ.a�h�B9�k�ŭ,�ڢ��G(��Y�1� ���!�/��Y'F���~�B�g7P��ނWb�rgI勃M�RRً>�g�G�ط��<u���a,з�t�hn{�Û\��,K��W(lR��v�R͖�QeO���밢_Ü|�@y����\��ԑ�L)2�_��)1��E�4��\������t9u+�̻;��x��A�y-��7�4�׺*e���u'; �֞I�~�e�_�CO�k�%�0�[�}APp�� ��7�4�7CI���x�Z��{5��W'�}�m#c�'I�/���?����>i�����v��V\��-�ƃ$������lG�NsS�d��Q��f�*퍊2ڐ��d$��)Z�{��ռ�����ġ�8Ի�T�#�K�߂FK��E��m���d"H���V~��G��.)w�)�=)�D��v��~�����k�㤯꫉Ȭ� ?�R�҉/�S�%3�a	c�/��q30�6�(���]�.r݄�����	���,;�f�'�v�W�w껓��*�ڦ�il��Y ������C��ϒ��9\dQ��8TX��J�I[7zB����ߧ#�lj)�A�M��q4�j9���R�)+�������]wD��
�O���6�9掟���$��7����!���F����{�'u�;�d� �E���ϙĜ��Cb3^&���SO�<Iq��*ͫ}ᴨ8ЫrH�=��k�	�7������rA����V:����ɎS�����	�l对E/35�N������;������(�*'Gc���o�yѥ;ш]�v�op��D��Ug���\�[*LyۍLJ��b~���dlTx5��t2.�)��ӎ:��ơ�]u٧�fZ��0с�b��̸�}�jz�]z�Z��9AGT=�Ij�ZDj�h#��SuC���|U��&w?;-4n���j�1�{4�,�C��ʵ}�)���H� w�V5�]�����1�o6Fr"��)<g�1%���~�!2Q7"��s���BR��p�����Kb�r�)8:�}�D<t@$R] �XQ$��N�6��/ҟ��d
�0�&��q�գ���lE�F����D~�ڟ�m�eD�� V���4��.\_k=&ˤ���_juK� ��>���|3�tC�
�h	�o`���ӯ����Ш*��$�d��ef�@.�\���0�}z�TTyJc9b���x'x��ĦC���s�{��X�ֿ�k=�ZJ֞Q�f@3*Y�޹����
˝8%����OH;bc���)@0?�=I���~t�_�O�ҹ�\�*xI����l�n57*bՂI��@�	�����	�ޑ75:$Cq��_溛�dϞ��~��Y*V��b9It�v�I/�f�'���Ė������Xjf4�\���F��)p��c�Q���sӨb�P���'������%L�,�Y��\�4�}M!'���JB��.[��#��&a�p�P2�^����e�ŧ7����H$��c�LC���
���qk�ByD.���D�N��5B�A����q�٢���i��3�N��u��	�񾩷wfWJݫ��O���9��Zgg4._%�I�M��+�żȂ��|zn���D˂۠�Ҧ�ART.E97�=W*�{��a����/���mX���bH�'��`ʲ�J�!�B�ܥ6�pVZ�y�SΣ��%kvN����]�莁��Ӡ=�J�)˸�-���&pFıfo`��(�AP�v)�o�彳���)��.�T�P�G<U�c L�N7oذ�u�@3��𰼻��2o�������ťv��y`.��fm�(��7�K4m�؛yC0~��*�\"um����|��_��g�Ĵk�z�������j���с��6gn�8�Jw�gkhr@^��.�ڹo��;���?���k#=�߉Zf�gf�	}
$�'�Oy�Ҡ}Xէ�Gl��6��O�@cf͔
������xp4�?������B-�:{i����C�E�O�� ц�W���<���=h�Z���h�+pj�G��hbJhcd`��$���֛A*ɱ�<�rX�P�զژ������:���aA��F�A�zrDi._w�T@����`^�������7	l#�ޘz<a�����߈U�>�ݙT��ԚF|�+T��jR�����Q6���^$�Lru<N��"�E�߭ߴ��)�y*E�]�G��{�4G���uh����M�k-��t����n���Ê�/Q�Z'��7"��~!��p�~��>x�XlxVHYEB    fa00     f50��[x�Z2S��\�&-,��QkX4I�K+��R��/[��+���w�l^dc��#I��$�𧏤׿��x��{���Aث
��cE,v,�U8
1�?I�K]b����N"���2��ȣ	�})_rF��c�fnS���%vKN�nˍC__���f�go�r��d�
�yT��+p[\YWd�z���/�V]�7jtl�2��U��H2,V�c$����*=���n����;#C�{�)���F��2p�Hr�:n{ݗX4gM ���R)&���2�i�f�ύ���N��f!���B��M�Tnmu�*�F��⶷fpƬB7
������[0��1��i��s�6&T �v���&e�
�(])��8�9����`��i�i��KW�Nl�5d��A��z���˩/�8+(�P�W�n������� ����7%��� $���{
=|3�[�~WӒ�.I�����x�+��{G���x~�� ֳ1�"%83nJ߭甓�����~ [����G*r�QU��X�p2��;�K���@� �Zg����ī�.؞���Y���,&��?�`�Ψmz��|R��~Y!u�����6M>�mL��<1�i̙����4����N�2�ὓ����6��2�(�D���ll#9�z�)����]?����kʝ�Sa����1u��e�!�NL�N�0�:YNT����Y�(�zf3c�'T��Iy�@ˋj�$�XI]7���%��В�i�;�
�ި/��U/�e��ꝸ�#�2�'x��ނ޺�Mf�Ek***F��m�p��'ݓdgw%����?��1P=��d��Z'�ރ����nȖ�����:i����7V)X��x?H���i����Dj�y�j����؈0d^/�H0��>Y�o ݾ�b�4�ho&gޞ���s?xVpT.�(���xD�T��"��zB��R���\>�h�a����o��^,�rIW�d���h-�ܟ}�!��+�g�Ts&D�Ip�{�s\Z����t�r_By�Sw#[�`�p�/��|��gv@,6��I����Q7fd��6N:#W�{��r[��-T��;9B;�����MC�����o����{��>�e���r��չ*��S���.��dvE��m���Ɯ�}�=^�Ԑj~���ʟz�������FM�7T�����[�Afhjg����M��D]5zg�c@A1R��K}�9M�������9>�AP������űy�	���aM$�ΚÍ�>-�̱{y�TƑ�ǩ������S����x��mk@�y�j3��
1O���M?iSij��]����ڈHr��3��r��Q��S����"�G)�Cs⏽�5�q���|L�P�ʅ��D���t���m$OV�HQ����\���y->�܍�T��s��$o�f 	�ic\Roj��WS�r]��iH�[�Z7A�-��訷��t�G�E{w�u����P��C���h5�N��r�Xۜ�r9�R휋��BcB7�\m~d���f�;�{C�e4νb��g��wfM:i�8&�|�Hl�j��M����a.�^_����{��;PTt�X��G�Z�( �Zoq�'��)t�f~�?ձ��U�sn����0���b�?���o�57e�ޫ4嬱R�ͪ��:y�.2�܈1-�ږN<Q�V,����|���`}$yJ���Edc;Q'SW��=e�G��]1����wv���	���x�q�څtva�n��������%b.O���v�\[��M
�q? {[!P�Ͼ-M�m7*�m:V� H9���@l�(׽Ή���wy����v�m�=Z{��_:��`?�F�A����W%�<u2���\+0�P��yF���/��翧��yT�q۸k�����3���?�p��-i�~Z�j�~lʘ�=��E�<��ӹ����ߎ�$[fj�2�a�&%]
&7-:C:�(MT�M��Ȧ�v�W.���H�d��l�ڃ�|x���s��Y�I\Ä�!!��v'�	㎪J1��k���9_�7O����O'��s��wV(��8��V�zE�[IG۹W1f��[�@#6U�F�w��ܟ����|�_���m	-��$G�I��0wg��^�5#]��C�l9�Ъ� ����W���<2A$���I�G�K�Y_���3��چ\l\��G-�]
S�b޳�U�KT�ֈHa�n���Q!������J�*�0A9.[O�>�g�m�\}���3)�-p���g���R�X��A�h\;�ggŌ���,�g����5���cĮ��h~�u9Q!��1P^^nUU�_QaYC9&����&�#�,����ڈ�@Ӯ�K���uB�p�y��Z	S`�[��%�.�D�*W���l���0��8 D����ET��8�c��ǧa�[���ǌ&���2���"����w�T�?�і�0]��[q
%�x�ݰ �aE��k�ޚ����wF���KI]���.��::L\䲩@�կ�'��H�`���{��|H^ n�g���P���5~�m\MM|��7#n �ԑ�wo�)� 6J��E;�����ղ����?�t����vEt�׳�	i�O�P���Dz��H�!Hdl��;�t)pz��{��vz�w��d���D���΋D�2(�y��_5��uY�W@�����m�����F�"LЉ]�$,+mg�b�p��YKڝP�!��T����Y	���΄��"���C�mS��=�{��|u�x5�t�A"��:>��1�}�A�&�hN.Sl4�<�Z�cj �䭝�Vw5O�-�����^|�<��t��uG��NJz����0X�@l�g߈�SQG
%|'��c���m
M,��#�G ���� Մ:q�Bi��T.֐��Ӄ��|.�F6ѥ,7�}ׄ�w�c�ZZB%F2�K��u��\�-,�9~����N%k7�`܇Sm��)J��?�$A��5�,e-\4T>��P��ρ�UD�8y�";�XHf��l�J1�z^���\ɕ�n�$Wû���t\3����,�8��)��Na�`��V-Ndً�n���L: ��eH[��5	�Z����ɡ���\��k�gq#F�j<a��+Roq.��d��Vaߏ�r䴳��|����[�A{�R)���AL">	�<A�5|ꚏ�@�  m�xv/ �m�d���"�+B��%J�6��C�3��I�R����̈S�)�+)(w��ƈ����4Q#�;bΆ�9<��Z��&�K�8��E���t�@����B]�ɉ
Ft�'6W�ߢ���F4V`�Nn��-'ۜ��)��/�^�Lv�Ǎ�%���|l����O_!��~�v�v�����A̶�I@K��b�,4�Yz���ԃ<G�ޏ�n���@C0>�`�0z60�KOK��Z.���1負�<~G��㏙3d
ڕ�7;�itM�+�B�6>�h���9�onO�h�����>��Rwo�9��L$9��@mHJ�)�b�+��ppYEP��C#�.�ݟ)<'Fg�c����T�Ht����� ����y9홅]bM�x/3؛��?�"���q!�MMEz����4~q'����Бo$�������J���h^#N2�?<�
Cr�,��7۲*�uٰ�����\u��E�b��Qc��P��k:�A<S�J�зD/f�4R�J,��^���M�g�\��"^wM��XK�F���n�c�19l�Kߨ�c������+�L 7��KCa�;���$�c�ƚ���U�N̜i�	�;�l;�N�0��;oޅ%:�E���OE����H���'��b�G��c �蔜#�e���gy��cA�KP��0�"����[T���8��XlxVHYEB    7273     560,�X@�/{�����|Wqw������<)d7'�#h���7�SәI�yW�FX�|��%YX��;�oAn'�/|9Y9zq��z;S�E:��1o)YAx��׻6��D�y��{C+p���� �Ѱ,�&�矂�'6��Q�m(�cB�ٽ��tn���\����f��0_����/�8Eyt*L=(�����`��I�'���~[,`���ْ��|/��lգy��C��Ѭ�Ey5�?�UfR����o�5����E+E��x�d ��(ς� ��� ^�&
U�Uv��M�XK;3k�2J�f!D�M�
�������>.�p	����;���A`P�j��愝!T䔅Hq�S�Z���i����M�3�:2��S��7h6�X	�TpV�Y�?ѥ�6����vX$�Y��hdL�p�e������D2k��"�8��.�K<(��$����BD�Jc�,�����n�Lݞ+k'᳆�a��n/�E!}�R�kM���Z}���p<>a���%�׶��|I/���.QT����ƴ�pS���;@��k�r�6�1����7q߯��.���)\ ��O%��G�t��У��Q�n,�u�τ	^�T/g4ߙ�id�E��m�o����;��|ցG��� Zlzj�q֩� �D�W�6�034�V��OA7����D�b���:GW'm�S���\q�.���xc��#�p��0���}X[�SG�|�e�>:8�}pT��e�: �P��*�R��ݢ��`�$�[�z�0/���3`���?
9���.H���I�'ɇ6.����X�q�����al�(,o�*
H�f��:*���NA˝���x)Y�yd��
#��Haٙ�QaU-�?i����ٶm{��qg�])ak1�3�Ы0���S�����Л�����F�}(�� ����J�Ng���a���ʽX�h�Y������-�2� ㉻6����?6R|�jr�M��QK�[$B�t��r���f��kb|�HD�P����+��f|���q}�O�����
�aU���R{��շQ'T�&�մy�����XTB�=3�-'P|�@:���'Q{i��i�<n@>��
5��0E&E^��j(@��P��p�#[�������������RQ�.j�|o�M2]������;�m&nA��LH6�J:ׂ���^7��6E��ێۗb�G&��y�T9B��*�ث�P������(h������&_"��@�<ˌ���^<p�a��/X��-~�;
5^�� ��L
� �kC�a�����#Ԉ7�|p���DX1����sy�@[�b�^��}�S0p�$��r�~\d.�hc�d��mZZ#)�*