XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��oT&D*<�>�I��]2t�'3�=�C��en��u[�<��el[1�i��q��*F[KG�;�H,2Q.׍_x�}4١u$C��k�Vqo�{8�Q]ŕw{£�K��U���r�<%N�ް�)���l��*���B�����2���f���a���S,&�+�|�i�>��"�M�3���*6"�����>F���D��+XIɽ�ӂ��X�_"RPAk�W�R�昕N��J����^z)Ԛ��}�	@�R�XJ�-�5�a�X���A�[���r����%ЧA��L�ʚq��&yLt^_��*���Qdk�A���\;AV��vz�	X͢^2�������ǉ�3�����3ۚ���;Ⱥ���!��������,t!�,s��+�o��*&��B��e+*����IHT�6{`�FޞJ[�ru�Vs>0���fk���Ɨ���z�H�=�}�hk�D{W�6H�"�'�Y��4@��	�������EH�{�|�l)�=�g��:#��ޓ��\=SR��N08�m9�2��Z��9�k�Љ�_�v�̟T9���v����u��j�>Q8^+)?�Ŭ�Z~�B�6�֠�obdQ?�1Cv~o�wr��5�r�x�Iܓ�n�6�����a4ɤV��̇��o�=�9�����_5�� � M�L�x�(X�ڮ��xQ�PFJ��Z�A�$�4R�o��f�)�w&]ͭ��ؘC\j�'|J�6�'�raa��`8���-eρ��o]����u6``ޞA��~XlxVHYEB    37dc     af0nP? �	TA�͛|C궺 &�I��Ri��<C��L�kvp�i9�M/�PW���hI/"S|������Ѥ���Z�?|��ر����4��9�]��L�æ0`7�2����%=�O|��Xt���f�,�;����՗܎!#^�@�zw;X���~��`q!��#^���j���׊� t$��gK�5�4�+�;=���N��cs��E���D�zv��F��v�E�?�����R���S��-�c�lgQi���J�ΥpH��nZ�߽��"�9�X>(!p�BD%�5����h\gշ����"��?X�dx�M��K����� ���
x�����s:�Hfb]�M������K���5x8�\�9�ֺ5{�[ %�/O|�V�Fq���>0����.�� �ey�m�7��r�Q].UxT���IW���G��t�x+����" 7

�����Mq`35���Yt��v�)�qՙ���/�]q/M�ef���z�e���L?&(����H︴��ٷRR7';�L�
��x�~X�R�4_�P?Rĝ<�U�U(���W?�y����V2A�9dY{���TZvb�&2���Mw}�c�HD|�
��{�F�ca�,U�����������Lҧ�|
[bו&�.}���1^?�)ǭ��TM��f���)����w	Z/�K|��L�f|n������(���~��Sh(&�r�;�NW�~���	����i/�|
��XO����f�?{��V[�	�]U%�W�B0�Ԟ��y��	)��Bu�N���Rqa��xrX�"�9&�q�c�z*'Y0��<D��"�b�O9����J�82)�)~��]��/�h@M�}PKBQ�4�^#�����S��䟊:.����}��E"�$�����b��g�^h�2���[���	v&�V7_e�a�D�c��F��]�%���$\lF����^�����̕>㊘�R��s_�����,O�C⇃S`�'�,;E_%U�f�)���N��5����W�N�WX��]l�<�a���������s�KrP��~o�	�rj�]H�Zp�}R���:h"��7Ό��AC�zVʤZ�.]�[_�ZF�P���?�I�������2H+5�:�1�u�ϣ�p�Ů��9�R���2�r\��+�E[���7'���pFO�X�p���ɮToq�����>��+^�=O(������0�l$��K½��y�(5 ��VF+)3�c3)������^m�*k�|G�R���tb<��{��n��|�1<�2�zV��g9��q��N{��B�[� Lz2����W���Bjw��bʂ�Y-��_x��9u���ĪհⲺ���+�ߦ
�\�\p�U���^��~��36�5M1O�I9޵xQi3�:"�a|�|TZ3�ׅj��΃��.��̝c����u?�� '�&x#���F��햨��6��:+�}aU�L������:&l>?IM��v���lzDr/�n���$���!��8]'��Wk�i�*�D���L[�Ẏ�bp_�0��|��Z�lm��)��]����m����x��E�	�4i}U:�ȇ<l��X��(ؕU��������'D'鸨������\:n!��jB�Ʈ���*�)��N���CR��7�e,И1pDΰа�;�u1�XaϥU���A+}I��fZU*\4j�.��L���`���8�yW��0Hz~��"��"4�́�	nJY�5T�΅6'Q�����b�#~3����-B�� �9��R��j}?�ε�oնZwp���#N�<g`FEX^�Z `C��=�Q��l�����o���4�����lТ�R��;ܳ8x��.5�V^�C�M��W�1��Q�r:lC�}�y w�.Ka$*�f��ٝ�L�ɱ_Fǧc
M�������^lg�E�� �����u�p�:a@]=G��H��z��
��7��<8y��g����+vn�*':Nj�|��Yo�����xhRѝ��0OU�����T��]�M����M�>\��B��P�����X�����K��dd<��Q�r*��X�b�ؑ9\(��h9w��K$�Ԓi[�=~%5�t.;p.��и��.�jC%�rA7��k��s��'#M�u�n)8�����@s&7/��!F�$�Az����@�I�)ӥ���+���u��}�8�Y��Љ��h��'V�E�pX��:�}�a����CrE�� s̍.��n����d�,z��Q���g�\.�-��Q
v��Ė��xB����9B^�P)����]�w{O�H���Щ�S�������v$���%{���Ƀ���*���� Rx3�2$�~<��a?�1��V�^�@����d�{�]���#�����B�#TA/.�(J���,��r~l4y�z��#3�6Oy<�s֟GS9iأ�M�9�����簣
ҫ~g�o}8�o�b%�\���ߪ.Vb����h�0�3�7�&rI��4���F�z@CD�S>"�c�F��K�6���K�ό陻����k�Y��e >Je�Z"쏧���WD�n0�H���ۑ/)6��"`����}Mfi'&��"yl5;K�l�#��zs��sa%����ځ4�~�p����N��;�>ͱ��}�!��HϤ��GQ�`�{;L��M�fO���ߛ�:CI" O��Юl��>b�k��AdO�}!F픈��q�
c����T�皶����w