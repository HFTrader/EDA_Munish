XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ij��V(�����W�]O;��YN���,>��F}��)h>��m�:[��~U�Q�\���X��L����_?9 �ӹ/�L�;y?b��b�7�͠ʹ�G9��p"�8��q�y�ʮ(�b3�&,�-��h�N�L_��<�}�v�	��oK�n� �|���5��vk��`$	_����L�����10���+����㇩�6x{�fF���d`W�Lf�	�2|���S�����m�I��d�`�"����U�`�C��1~�2h=<Ll��:�D `SS׸;��E�7C	��Ջ�N%7�Q���)W�ą����r8=��� pB�J��<�8�D��k�H �"b��^���v��V��K������)2A�;~Z6OU���tx���m�a�~[$_hg%Mdf"�@C�ޡ6����S����G�:N��Ov��c���a>��S��c��7�WIs���eX�f��ΛW5�;������I�`-�P�+�
r�oRf��%/����)��L|MJ���pj겢�>��T�PZZ�n~/�a�l�;�-Yn����� o����w<i�6}j{�����򬔷;�����ķ��)E���;�U�ջl�М�|#f�CF�\��[TI�4i	p���,��`���� |���%A��w!Q��Gn�e?����?{�;�[�=�e�E3dW�77�[ļ���ѐ)e3J�������I��(����EU�cg;�5��!jy}�v�2Gv��t8дM�˄so�MXlxVHYEB    6534    1400��ר�e7�s����
�"�bj�*-p=�v��b�|�<p�e���%_�f��7�)`�R��6�']�����6�,yum�I����������9��;�w�����N�tXdC�(zd/�C[#�:a�Tۘ�����+ɑ��� H>�>k���¿�_�i"�Ҏr� S|��Y�����}��L�$��D�����:!S�qϕlb*٦�9	�(og���Y�\��v�J�1�_�\�N�zj�$H��á��m���堾�F������ZK�1�]��$�>�Ͻ֭k�#��1WgT	�B��a�m�,)��'�Į
{�Q��f�l�f��Nci��O,��VjX`��^��PL$�ӽ�t�?Z�Lm���es����~jdsX(-��\/	��ʜ!���J���:��ʂ��D	���_y�|����:}�`���U'�ڎSB&�]�ٚ^ �[�K�:ڲs�%����2Ģ��������2�)�>P��T�!���1�^^1IӅ=R���.�@P���|�[�g���m�f�������g���_��	"䌛�y��f�x���{�!�(.Ɨ�"+�X��,廴<On )��W�dΟ������ea������UM�Ho�����"��1֔`��Ȼ�:��Ty`/ְ}z���A���r�ƹ"�J�}ND	\#?�g>AF��g����,-n�Zo]���S��g��<��^���E��1����Z��Z�{�pU|���J�Fwd�Ԩ7;i��jo�?�^M�L�����K�������k>
@���|f�k���m1˧�*񤞂�ňY�U��/]-n&0a���w��D�]����lIwŀ�k�V~��m���N@����e��)-\�w���g�e��H�y��W�#���N��"ߦ�*Ȟ�;&�P\����j.j� z�{B��0���~�j��83-5��`kC�!̛��Q�
�"U79�� P$�Ús��Y�ɾ'�M/	��;����p��s��3r�8�M�DG�.#\jy܂��X��٩ց����T�I��&~wj���L���f- Չz�-mb�r5��k�	-6��@z�P1�rL��D}��E���$#sf�����d`�e+�%�1�
n�n��T�Tʑy5�^W�><�����ӹ�y�e$�٣	�\:�/K�ʦ��_J��r���@�uf��+w�$>�m&� �]+�]�P��	��ex6�!&_'!1Jn� ���^��� �p�0��@������Fωʖ�����޻TC�3�|ڽIL!02=�?au`��sQٻ�^���8$ �j�e�;}�D�#F���ㅧ;��Zgv��q0F'~ڌ���gM�����i�g������OA����h�.;���׎;��J$�*(��8�z}d?'�_��|X�F��o��x�5H-�9I��>2�-}_]MN��0��/�
VW�iz�7DI�@G��$|��b��dF.=ږ=����P�.�󣌈K�@��Pb5M��^wW.����G����o$�Z���}l�*B�PJ�����с%P4Y�h��S3h{E�:��A@��k�FWT </��xr�D�{&q�Lɍ�~ͭD��{l`)/L��g��C�)��s����$���������f�!���m�*2��ʬi�����������u��S�:��*8��X���B�v���c+�����Oe�a-.>ˈx��{�Y��k)S&������ɟÝT�{��q2�4~u���~fa�\�7+��g�Y�YI�#=��h[�>��~G3���-z$<�|�!����؅���`�Q*� l���]j�����<���x�z�x�bcF�^�@��]�ځ����=f����p������,Y�l�HgIї��<�@�8dZ'r6	� �F��aG�� I���Gj�|\�ﱵ.�(�]���\%�'e�Yh�>C�6�bƊ�c�X��G��o�G�ɱd�԰ބ=�"�
��ci����J{~{i����9��B5�HMD(�v$�!�x�f�H�1j��(�~����G�}o9�%n�u�1���$�I��C�E��5���it>k��~�x�r`�s�:��>P�C��<�A����)�7��
s#(u��=���;0Ԭ,18�0fR4�%��#�;�zt;qv��(�$GX��J8�4��/�֩L�G�P�M����I�a�v�ν��q��B�S&��\�f��u?�Z��$P�bU��T�/KuW᫛wu�T�w�_ja5P	Ec��%�Pb�/	��p�AX�-4c�H=We���:pAc����\�9��P�qH�q� Q��K$SU��^kF���M�0>��31RW�1p+�©Z.�����τ���#���A�li��3�=ࣷ��gHW�hB
����ζ>`!�o�|�֮�[�Q*I�p��N�4�C�@������\۾��4����8�n��%���U��R�6�0�lx�rl�b�~��.%� c\dI�-��"��Ș9�B��j'�%��;�+{�'�7�Q�k�_ �k	��bckq��M2I�=��A�\hO�״Ŭ��8o��m����x!��h��R�3��/�`a�)��R͚MSC�*x>kt�f,�������ƽ�{,�~�伔eс0Z�:%�^�ٸ��F�`S#8 a����^��o��ҙ�g0����V{P��B'���}ez�3��LB�C��Pk�_^�J$��T��^AupIXϐ���bs��xȜJ� �,�q�<iB�D2JJ����pi|�|,J�.�rӢ�,�t� P ���a�3^2&5���u�ǿ�Xy;^~xH���6r:#�\30(��V��N��fM9^a�k?�`s�_��~-sk���e<�;iRr��и��67���%ѷ�1�J:�w%>L���N�wq�D���]�rU2��ۼE�0}�fm���{��U�n��Lj x�4���n��ScW�bH��4] +�}mI�/��#�FS����*!j6�� {�Po	�cSJ�%S'S:������M�<BS��
�	���2^F)-�L�5<j����jF-â�O5��.g�ﭠ`�7����}u�>N0�2�3苽@ů���A�:��Npt��p�'9����W~H.����1;��T��i�I�:ڭ�.�����e�ke�t/��|��室{;J��4��֬U���nW�)���������?��5�#��_ A�	9V�l��y�,9Uf��ﬔ}:t��	A�[HUeݬ�P�"��+�D��������-/�Q`B�����5�����K���[���V�F@��,���J��u˾�~B�,�iNC99N�MHҰf��N&ˤ��Z3��,yw��jCo�"Vk�Z��#��LF!sߋ�S�σLW,��ѕؒѕ�>m��m�"
�!�P���E���V��H�k��������9c-�,��l���B&�3L)�'�����1�n�;����Oi�w�g� ��N�w��
���SJL\S���0��̫ˁ!4LTT�l�|���8D[
Ӝ���g�M�RڿCuU[����S�#���u%#Z��N44���s�{��G�lf`�*/C֒v��mG�Y� �^p��.p�2��e��AbXk�l:+�6��_2��B	���`S/rU&AfA�0��R,�^�51��h��ݷ�AJ�͓]��Pf�e3��b����M��3�������|9�U�@zj��*#��q�MXXA�� ��H�V�����Z^A�8�ݸ��ja�i��\O>����Dp�Ya+�aG�����f��2�ر���ԔY.�X�hF���S��.��r�D�v~��>�㍭*		SdXf�Za�+���E���`���+y�r֚�S-'Ϛ�W�W/����#�=S���.���s�PH���ܐ=��&�4}f���|�4v��`c�>v�]�t��[�'�ǧ�����"g]m�3.�x�j�	F#�%�U�"�++M��z�Z΂�������_�ơ�h�?�j-�u��5�
���|��,�+C�!�N���:>����,�Ϣ��;��?iD ����������������'�� J��ߝ�5o��4^���\�髬��x������ņ�b#����c�A'ԹM�w�/��Y���Ǽ� ����n�h�;{'�3Wf�R�E<�}c�VZ�[�Gz�V����i���i��������ր}�^��]��g�<xu��w!�y�$I�
�p������3y�)�UO"2�����L&��fJ��ah:5A�Ǻm	����rx���=��aUDZh�� ����|��O6�}U�3�c�p׏y�r�x�`~T�Esu$����J�8��
��C ����(�#=�r�Y�T�v;7���ޗf'���y�5�=\}�l�UֲZe{ܺNw���U9g����(�6V�1��6�G�Ѝ5���.��¿x轊"�l��8t59y1�o�1���T|cj_Φ�"�.5:��sK�flo�F�3���3�vz��)�����P!ʶ��U��B���l�/�X�cO�em8���ө��LñU!����7��x�B�(��ٚ����i�,�t��2f�A�0y0����+չ�B
�2\�-a���/)*!����yͤP��C�4n�G~E�����?�0���X��9�1o����.�E��>a���A��%Y�c�#�����K��G�I���sP�H����M�@�v5ZT�t^3�Ew|�֜ �DU��O0IR,�C�%@@��f�m�%���)2M�Q���%���C�D"ھ�X���W-ԋ�do��͓gc����C�}����D���;'6�Ar~\pst$�(�v$�=s��N/ T�S�WZ�}G%.Kc���]��F��z�>�F�a$X��_�����q�r��,T<�b�(�1����'���x�Ms�uT��X���[u��_�W5`�4�ۊ0��ז�B��d
D��P�C��|��}�\�"�������Ξ��~�w����B�E�F�7&�{��U��L
g�@��jJQ�S���