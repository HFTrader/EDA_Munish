XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Q�ȁ�ݡ�CA5_=�V�����C�i���1��&�VBD�6VAq�'������� ����Q����]�dٿV�_+�|'m
�T�>��7�+7X&��{��s�z�ig�T�=��x�>���ϫ�9�e�Pr�5�P2<��H���@"�]�X���M���Õ9U{ ��ڼHm�̙�i������{��D��m@�����<(���}Q�e{�ߠ_�0�" ����*�m����k�2���]���LB������!M=�_U~&~etrk!@pO:)��t���a�vH��c��b���ɿD��?~@snK���w�uU
��-�C��GV�AzEʙ\��
�ٸ�e���,z�ab�xC^ي��'�.ĿNAE�H�#�'H�%lP�Z�r��n-N��_��1`�qi!���ޖ�����<��T�e��@�#ݗ��k�94�
H�"fq`;ɩ2�;��NHWAO�;#�1vׄ�7}� My	t:َ����۴EGŦ���/� P�5~����������!R���G��?{�Ydz��#e�cn��a\� Z����/h�����z|m�k`�uW ��
�c���*���c�>�T��` t�E�+���h�Vs$<V��5�vC?��&]�B�\��bG�� =V�k�$i^�8q��!��ȥ���絽���^fr/"?�E����s�:�u4q���pa&�;C"��}�������L< ��=X����XQ��z�CK߀�Ic#�w��s�P��v���Gx�Ҧ��XlxVHYEB    3da6     fb0Z+"��s�p�~x�iȐ����g�y8��ښ��f��9o�2�*�.5Y+, U<I�"���̿��p�%GBH�X>��`϶!q�M�|tب\��em=C�aJ�9�&�G����H�.���B�kmg�O�@�tF+�������*ݽ�`��w$ӯͬ)5K>��<f�^�;
7A�tm��DZ��lKb���߽"�H�O�6��^pC�f�_���bLH5��]��v̪B��샳��ݪ����k�+�W���	��/C������ƅ���DiC��6�wz&Xl��ҁ8��IB���|o�$E�ˁ��^-�Q>+j��r��G��/�~r���iJ#��a��q�Mj��t��F�/���ۚ�<���⒎%7!Y�4���fuL@S�;���RqD�Է2�`)�@�8�@w�a0?�����A1���ݭ���Qt){N�5&�8!'��#�5��yY��&6�Oo�9��d�^��q�|��,9g2]�G��5÷v�׆8�"2A�_2EO_��^w��1����0���/&2�"�o;��R�bpݷ�:���lM�f�,eF������j�[`TB�F�Hԉ�1�B��x/5ۍn��	l�c��g?�:�~�d'�e)t���2>�A2�շ���.!U$Ouyv�C˄��R�}\T���_{Ҵ����W<F�����B�@H)o�[������11��B3�����?��۵��T8�x��$���:+I���dsj~��^��\�Igb��'nb�Y치���?2t��9'U�j�����4#�2ڤ̵�>u��SK����%p�V�O)�h�	��ݚr��-?�P[�y��a�����0��+X���1&i^P\�����L�Y^}#g�. G)�����k�������P��;�2
i�-Iv�]ޓ�����X:�m���x�OpSݝ>��Bb���"�+���sT�g
�ED�M~MS<�H^g�����)n93�����妟@�%,�*G9���cf��a���hyԼ��d����d>�cV�@߿MF�Զ��IY��[�c�6�zE!���)=�_hU�5e����w�ٱ�`�32:���WI��ߋ�eq5F������8y?�'7���T�ӘC�s�4PGaݓ�����ݡ���WM����se�ֱwE�T	؀t޳�1/Ni��uf"�$�N�8�s%���K\�ty�� ���!�xD��׵��sC�T�"cxvV9;D�않8q�8��Ue
�ﺍ�o)Ja�j[��j6�1��K�:n���& r�q������%�C��{���W��]p<������7���\���bw��ts4���Y�Sl<y�XJ������N�"����ʕn��gs�R�2��/`��a�4|�$�����s<���˔�±A;� D�%�5�d��n��l ���	FMӲ�v��oM�۶N��`�P5��v�	��!�[d�}֙N�l��_�>���|�৙t1o�J��U*���lq�.�U*�A��f<���	J���ѫ׈��&�z��d϶5Lk��5�PT�c}H��FM��kٔ5�X��Q��(tT9�>90u�Zh�f������ds�<ov+0�:0Q��b�P���%Q�t�a��C�{G3�C:@�g��S4��^se����4(q��@�L|<ۇj���pT��U��Y �5{�^�0�&N��OB
A>�����		d�������ϸ�SC��U� u����[�d�Z~C��E�4-��C������9��`��x�"��'5�OG�H�u��X�E�!7h��GFk�	�`��@�u?V`;�w�@ٞ�=�d�&�@��Kf��;���ˡ	CšK�#`�!tfݭ�����~�n��lAi�`x~Q�n��[*�U�[��Y��7f�a�j[�72@�n�|)��j��3͖pz��ĉG;E�]��>T�gMv�v�/ל�h�x�f�~���,�^/�AWC������8}�H��儡�RY ��Še\̵zד�ق�T�K����+��T�Q2�"��V^fA��x�"<��ZZR��Չa�H���� �������z�m\wLU�,4~�ӑ�DK��=�#�烣��b�O����¿�j[
~i��~�d�CE- �-��?��5����.��P��e�\��;1 x���O�L�� N@�6�|�ʚ3L6�8�[��E`y�L~�i�^?;��:�<҈� 
Li��b��+�uS��=@F�}���Ϸ�\V���b��������SkTO����<*P�)����謵�7`S��Wp����ZN����I���֢��}���Ţ�� �G�_��\�
A�����3NW��.�M�JR�dN\�JP�p�c\9��i�1T�*YI�J U�ҕ����O ��\�����ˡŚt�c�t����@/1��M��V���}��U��d�;�"�t���X��6wO�@�H'3^��z�L��Q��]�J�-ۄ�(�D<϶}����SMd'?/���9�k�=nVW9x`������/�Y���t�V��/CU=��C��`:�0ö0�T��o�����"��)��b䫚���GU]�4#q�i�����[O��Nm�"��_�߳�ҮOUf�}d�W� ��aki���mr,P?��sG����61���	�t��Q��w����(�ɉ*pe��o�h��|��WtƜ��s�tAt�f\�="�}�Ԫ�8�e�@��{��?O>:9��o�)�y�]&q�;��,�`EN�2�c��	��� �`���즓_%�;s"8����f�R@�ͭl^�60HP�~:��=Xu)6�" a%eS���Fl<��p0FCO
����-
OcF�r�\[څ��}�f?E&2-L�-�-]h���K�;�ٵ��Q�gLq�9o����.m�|�Z٘z�]�1��-�����k΅�����` -�Ud�Vw�[�dkl��Yx��B0��@�A>���+7r�(��q����ѡl+�OB��B�+�J�(�CͬI� ��h4�M�LG8��ϑjl��#-��4������u��h���������#~9�,lĨ�:IWt�
�k�8%W=Y��2m�Q�.A?+>0���gʺW�?�l+a:)��P���a�J���c�p�%�w؛D>�=��be�m���v�H� ��k@�+��B��d���T&F��E��U��A���
526�7]z�G�~�I !����� ��:.��crb/g��Ssf�k��^�]��s_�p���Iwi7���8�d=]��$�Ո��8�P�-���:���t���� �{ҫ�T��[ϯ?ݖx'�%g$��a~�DA��J�!PST�������V�=��t��_&nw�0Cߐ�dh@����$b�B�nw!D�cT���-�:}Myv��Ս�#��:��~�ʎe<{�^%r��`��E(��b��1G�j_�夆�)�ߎLY�(���
�[_�:>��<��~y]�� zٱE��d9\���'B�L$��)�H�/Y ��?�=k�P�܇�4���j�:�?���X���k�╠���|o	ȼ�n^�����?�t� ��ǈ��x�f�o^��X�Y���.-[�m�	���5�٨mG��b	-M�� »�?13���:w���^����c\]�y�oi�`�:����[�8��k�d�HN�ɐ7Uރv(�T��e!ۘ��6P�vzm3`ۡ�TO杺������]'s�0A��U��˝�ٓCf֋{c�1�&���\��KX��{�[2��yh^&��=�(_���
`v�Qmk2v�qZ��M8y�u1�?�����m�-����͏�Y1�����Blq�Lq�������<|��ְC�Ǘ_�̩RJ�v��<`��[f,�ט�Nٌ���k�M����}i� k���!��H��&��������fx9