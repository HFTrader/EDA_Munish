XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s�����f|<{���{7��P��܀t��[�7��T��svJ<��c�<� s�o��O�`F4�����\}B�'�i��y�:��α2pyB�ܖh�&�+Ux��u2�;Uo��,�=�}-�x:{ |h{>:���w�p�b�S;{�w��E1��@��������m�\��'�y��%�Fz���.�����
(uo�s�i�I�#�O��������'�&���L����&�����}W_�@ŋf�I�D�n�lΜ�
�nS�3�i�"[��7�M��E����C
/��T�4�*��(��:�;;Wz���[3ؓo0o�� Ԃ"F{[p���9B((�@߬{��l6���'�wS�����}к�W��U42��rIo7�fL����1��D��'�J\�j_�^a��X0Kbh�s��R��HnԘF����d���'h
	��$�- t�7�ې�"3�k��Nm�p�&1R����\�n�ڌW?�M'@gEb�)��O�[��Atd��vnî(�Ԅ7o�@d��;�����Zu^����)�3�S����k~�#ՈCL�K|a�JJ�#Ɩx��:��[~#�9.��0n��nv��cV�Ô�᳙�Y���`����?c�k4��_���Z٨f�g�#����8��S�U9���*2��n8T�? ������%�N�@���.c��UB���.���ew�x��%��l� �A�����)sS$U���wU2�]0�d+�  ���Z�B��y��H^�ǫXlxVHYEB    d7bc    22e0�Q:�Dc�6����Q�,��Ϲ� �ʐ �^��
��s #�|)W�`����'ػh��<�[�����s�wZ�W���d��.)7��AA�B��?x�8�Up��f�Sj/=�?q�����-�E�����,��~�ۊ����A�ת{��`h�wh����'Pb�e6��Y}/����Ε5�eH��	�����@4g*5��ø�Ǹ�d�:�������ص�&a������vb^@�W��R��^�E6�8Ѷ:��~����)XԺY�w�c���p�mFs�V�d\#�0����1�SLϘ�J9[��..�|�}���	�<H/��S��N"/�ۖR��c�����D�"ϓ <95ꥵ�ԥ��8��W�[1C�Lo ^��l�Z��En��9%�[�y�D���A���*�s��֖��n��Y�>�/����Z��I@�%<����p�l
�'�G���1��!��~!�*�-6�u�����j�����z�1���b�Dx^��&���>�.�l;�JpHe��E��r�~���?K;,�I!�X�BƐa�h~��0W�1�P��A�,嵇,/r�u��b�؊46εfڧv��n\���������lv�����]�4=�p�nܗ�p�[�{�T�[���#ٝ�;d�,��AQ݈C�������?ˡϠĺ���#��`Y:��l�󸧠s�S�t�|�@�_�T��J7o�PT���������� /��~�˿��eO�af8��0H�A}.qcs;�WRS
WF�r��qT��uD��K�{�y��{��Y���ym���p����	+Y��+�v�����~�R�K�6�d�ij_�۞��\֝���7AR��S�g�5;F��q��s�n%��n��[�[V�yU�����w�4|�T,28��AɔS@+��*��5�[hBED(���j�@���dl�����zP��%F����plio�Un�5n}���3��2M��q��͵,�)X�}��d�H�s�#~��q�ٱ ���̫�a�^勁�y*E�Č��ɡ	Gz�"��ߙ��/���	���Rwq�r��,�-Ʌ%Kj�b�dW�����g���n��a�\׌7��1X��(����P_���z#����]�1w�c��AScnm|�T������W�i0��.φ�ے�R{��w��x�?��=T�`#�3I�Կ�y�U���Å�i��8�n�"�����C��Pǆ�3
Re���������8P{+��x ���ǃ���/&ZU�B.��)�F������*[��g*�����ړ[�]-��}� ~��r���[L2��V��)\��9���7�Iޏ���`f��pC�B��HŪ���D%'�f�ߵh����:���x���,` B���		r�R7�c�^@ ��rw>���ۏ��!8P7J�#\T�]M&I��qr����"���՜R���xO��D�%��y}�z9�2 >f	@�vKfpQ����αsxM%Ʊ�f-din*�hcƪҖ��y1+���noG�BrY=�����4���~�EWS�[��X�:S�1�!o/�y���ooj�'c�NP��(CUk���-� ��Z���e�ɜXBX���a��'�s@.���9���]��M��qmL�?8��.��z��3�%H�T.8PU��[_�x���c#3e!����Uv�I��˸�j`)��		ߙ�7����I�d���S��rK�\R����A�FW��%���DhE~�0�Y*�f�LF �CN�� %��8� ��z��X��Q�K-�\�A�+��K8䲗�Fҥ�Oo�]�\p8�VAC�`������L$+��qo܀J[�֏�t��@��Ŷ`\ԍ���}V�$�;�?Ģ�o�b��[20q%W��hwL�H ��Ï�O��hמ�Wr�G
��z���UE����s�K{��x�ob��Nck=$KjG�S��B��ol%�+.pm� :�6��n���pW+�3nF��Js�<A�C��Z������d��}�����vǞ P��X���\���� �`Tmit�ޮ|���#�i����f�a�����O�Q�����&E���7*/���	F�;�2�mC������e�GP����HP;3�.���z.�5K�>R�L��3��4gv�n��ՀĠ�ek�}Ph꽋w��@@C?q*�Ё^���c����d�xg��=V�aX��{P�"��w��/�5|�>Ȩ1�#���>�T�i[��K����'�1Yd�$f���m��ֆ��������*��V	����m�,_�pi��`ͼP56r�{��ʡ�f>���Fy͚c�>SN�FY�k|� t�і��V�����[��0ĝD����;�j�KI��\���FRx��z�!$ܥI��k%[�|��Bc���U�E�Ք�K�����j>��>��a.y>��e��	�c�F�-5m	�����G7�40�"K�i�$��@�����*�W)���ѽG��5�l�x�G���]��]l�Y���b�)�IT�L�F�K��M*���q����ϻCVcI�[�-�W/a��
H�X����9�����Kv{�]�؂��
�$a�z��b�s4��+�G��$K��5�+"�����>Z|M�P��1�Pc$Zر'.�h$�z��G�¤�dPl����]�6���dӅ@.a�e�h�""��� +v�8)� ��^86�����D`i�'�L��"�i,⿅n
���<�����e�s��ِ�ULK8���#�6����H,��^�p�j�`92���N.*��RY�W�q����&�5"�#�K!��Ǆ��c�!(ָ���D2��%���Dd#�Cʋ�L���D�u;���o��4)&P�^�XY��`����=�o�Q�l��u4�W-�t��Y[!ӡ��hk�B�T�<K ��NHY���Z�x��ctVy��^���(�/���#�4ڊB�Df��PQ6%��\�6��
�tT��Z�%��۝qi������"ow\��0��S�X�� ��r����̥V�vV��P�r�����]��FT��r�w����2�SK� �<{�H�um�~\�E�|Y�8E�\:�ݴ���|$��`��^�	������LQu4���x��"������C�'�Iا��;�?��{�Z�+��!|����ߓ@�V��g�#T<GO�*��uWO�����1�7>�B�?�i�p��x������<�V������\H��z��]��b��p���,�x�lȑѫ7�rS{�9F�~\��k?p��g�D���5w;Z#	�c��@v�&��Nm�r8��٘/�����c���,�U�T3��k�cѷ֎@�)��pyç����ꅡH��_��a!%����7i�Ó��������&�����#mq�U[�F�ERC�;���ߕ"ޤ��U�t������bԒ�H� /U��d�a9{u����{�'���������*�<�}(��R!�뙲X��g��[�.$3�+4��솋����y������w9�T>���X,�o�y��U&���Ɯ�"������C3����$��X�T�e�~��"�"��	�Z!Q�~{h�K_r�
�N�p$�Ά���DX�P�T%�ވq�8�$ZD��c�I�ח4�ء�g������f�X��rݜғ��X3P�R��٧X��Qm �r�S;2�$O�N��_� �[���F�=�\&
��ڪ'�Mv��Ѓ\�İ)o�LF�եP��9�'���r��u��J!.M�����'6�n������iF�ҸV�� �.Dr��� #��%��pZW���1�3��_0u�祂�� \� c�v�Y��'���a������C@A���B=�DMj�э���t��N\I��@�������.�e���P�rq�p�^IB��W��������\D�ܟ��.�/{m챵l����\.~P�W�tZ��E\�{~�x����Ԇ�����6}H�� 5�hu.e�
uI����+Y�Y����L4����n�ޕH(:���d"�x�y[�X�p<Lks��N{׎B4*�R��.��iW�L�&�cu�W*�#�s	9Y��d��x~��P��Z6 v�dg� *��"��IEv6��	��6sˁ����YW�k��`P����E��ǂ/S(��@�ƹ���Z5P�@���j&p�*¼�[20\'S�>;���{v��'��4���n23�;�U��ņ�Y�B�'g��}L�(ĠF�'��q��{=�?����q�*h�N�Eh�}&Z��%�/�W��!
Y懠���d
ؽiHU�u�d_h]��8�0������R���۾�U�5��&�)���n%f3]�Nl�/Ց�):��H���6�s�z������l%��*�=���\������t>�u��dd�7�BR;�[7�P#̇CE��3
R��d�
��^�d�+�3�p����l�(�u�^r?��"/��I��T/|�EB1/�X?���cdQϏ=s�W�M9��}C���FRUV:P�@�t����~��1�~�Lk����>�И�EE@҅a�;_�N1�#���)�䑄��u�S4���a����w�/��B)��U��#�5p�.DՀ��J��Q���ڼLe�E:g2�������J�m5i���^��i�hbcU��*a�Z���5���(���OQE��J#	cRP �n��jId�_y.(c�3Z�+Sex����$�XB�Qk�y��|b�̿\N_�I~���S�#z9O|s����Cr��~FV�mtoz���ynkG_<~�q5uS��Lٸ�!�hJ��Y�Ni�w-�" ��J�j�.>L��z:�8�v��huD����]�m��\��2�!<��AzCy�x�K���*D��4-�0�����h����n`7(��lr)8�յ-
`]�[�bz.u5WWx�U�!�.dh!��l�E��6ŵCY=(�y���R�Q]��;<�8����y���
����9ւ�ؤ�AC�4`\�;��wZ�?$�9Rhv;�Ɣ���$��[��}f�v8UT,͌����3!#Kq�q����C�&���X2��e��jp����$9�ε�k;�x?7B�z�~��4�fg��":�#{K̙Q�pSwT�m�^Q�6�;8�lt�@OG��/}�����J/v}6%Ҹ
���one]c�Z��j�-U %��������3�7 ��b�Br&8�DM��؝jW��yǊ��R���gL��ﺠf�j^Kx��M=c*;&��n����Ns��Γ%��7�;ܗ�St�zF4�%�Ц���<is�X���i�l��R����2hX��"�B����y�w���H�4�_�IسF�T�_���y �9��\��XJ�P�s�n���v���I�,���%=B�Fh�N����{��r0�ՠ���] �*�'I�4��6���Raw*M)��2/�YH�^`n5��00΅��K=ߧw�AR�B�-�ޥ�u븹Y(�5�	|[6A���L��	��m�d[�4�a<JM�mktA��BS3Q]�(�@�Dh�Xz� ?�#`�����H֧ױ,�m�$���WQ�*��kt���+R}��
])?� јd�]��	�/�@�����Bu�ִ�g�8�#ô���������kn��8߃��*����<c����S" �qN��S�YO�ny�c�Y�0���TNmVY+��7�4�.~X����4���M�a"^&�r��{��v��i� ��oW�>�|�D*{X3�:���0������ք�Aw��%�w��]�k�����s�r!�X���K���W��Ϝ��!���e`�� ����G�r�CH�AeU�l�F�}ס!��e�ofM�����l��n��q��ag��V �]	1i[�Ī^kҺ��B���UC>=k�y�
�2ܝ#�+�_�sp�*�g�Q�HY�n�!+�WzDdq"���We%%$G�����W��X���D�=ݙ�R|��_ʃ]�BO��w�\�Ɲy���_=cC��M[���6�@Y?1��$X�@��7B$q1��$8�Ya���Lqe�53�������jV5ƏP���l�?��x�,���8����8����e\��+�1���{b�%�n�{0)��¿��l�L�w�kft����й���}us,�*��pg�v䦂��1�Co-B�𕞫O���	0&�^�w��8OX@l�D q�,�IF�Մ�?�c4�yw��k�_��{��� h�'�wh�9(+]"�姒��4�$@TE�9C���߇�R!}lLL
	ix��z�S�\9T;��k�Ӄ��ր0+��L�$�|�|�n��&Q�z��o�������(B�{�Ueb<:Y�h n{����L�r��Lص�-��
fԫ^�}�vO+ܓ&�W4'��>�'J
5s��E��_�~l�\}�������%S��r��J�B���Ly	W�%�����$H%+��{���]\���B�=��9�6�c�D���+#N�W�Q����{�"�h�u^�/qEG�IOo�a�*Zv٤ �8d+BL������wc]���0��1LZRT�Y�K��'�
".0�t��F^b���� \Yw%Z��̀�c�"�\�,9��ߍ�M�6�����,�!H���|1«���!}7ɣ |�d����֎g�`�C�G�G�4��K�FF��k�E��ӡ>�Mީ�c�׷���X�j	a��J��^�,ɤ#�i[��l��O���O��q�M�?A�a`쏻��<�3`Q��j�1�`W!RD^��f���.^��!�(�-y~q_���|͎�`�h�2�]+N۲E��¯��#+6�}���A)�p� vwTd�%P�mmA�
f��>��PY�x�`��a��%f���|�u�]����Bx�3���A���Z��g�d���F�f�Ⱦ�!Eҿ)m	b�T�*�E�;GA�a�¯��޸&'1	1'�ˉLj�������9Ms�
~��c� �uv
�N�������غ�eJ�+Ѧ4���9ϻe�'���%N�X�����(�0w�~�0K;@�%"rr��.�1Qo�u���(S&����9(n�"�o����\󘳲>�\�Oj�q�g[�Y"�<KJ�fMCY�N��+#���"q_�1��o�Ƹ���Y��2��mDw�[�l4c�;^�|f-^+���0^��_����
���/��>)��*�<h������-��m���vA��y�2���9�8%�v�!�� �Ӄ(Y2���+X����Vu����o|��(h��d�|L�ї�XcÒeT��ܠ\s�`���Z+��`���T|?����>\��b�F5��� �KfT���~W���})�vs����8�:��2;vH	J?�93��M	��b�@X�-�e)�������A��]�����!�@@�t:C���3��6��حle�d��-�OP�2��҂���W<7�rKaD �OB�9���'UUPr�QͤsOI��KWƚT��Q�|�O�_h�["���7�OU�`��<fZ�2Y�lu��n��c>�"%��W}q�|70S5�$�6�Gs��q�J�Y�*A��I��ɣd��q��oi��/!b�����u\�^�R�2�إ�n�r��e�ź����TR��1�dY�0��t/i��u�0��גL�b\��4B�~���x�|:X�4;�Ԉ���(I}/���V�i�M�?��c�Zck�2����qI���:N|i�#!'g_'�hb�ߒ 6L���<�ȧ�7��ݱx'q��ȹ5ʬ�Y����Bc��J9Ş��1mE���7^�������p�UI����ق�Z)�\���>���#e���+A}K���˔-;^\�╢{�k�֕��.5c�p���G^_d��(E1�4�.%58��H��xB"e�|pv7d�6��.���{o�·S�Ѳ�D���ܻz��_64r������OS�Ha�2��v�Y^`�"{W�!�=zF��:�'��� N
�˺Cu��zǙ���m�J�@1�s9%J�Qv�B瞥�Y��p���k=I��y�)|C~����t�3�`6��b?V�g#�Z3��V�Q���\"3���,���ۺ##�mMua��8اp��?i�!A}�y`�HiF��0!��7�8��R�z�Z�eKZ?�=Ҽ��΅���>����6�<�\��Z.:�Z�QmX[ɟ�Wb�F�h��]'��ּJ�3�7�mˈr�c�py�eǡGլ�����I t�;�u��LM	��v��C�^��k<Nr��E��"]w��H�>����E�h�6�R���)����,1�q�b�Y�
��������z��!�]�$���]�FK��))�ʞ�Ji*p�ݕ���Ӵv��:���;=�� I����X��#})�UCg���_��M��DW8�Q҃ȸ4��D��}4�x�le�H���6�0��?�*�
��^]!ܽ�T�~�wt��M�E�5#.Q쿛4(T�fee ��˪[��>H x�*�[f&s"�[,���W��@} �f�ums_Z���4���z}n�/:�!9G`�ΰD�U�!��j/����O2�?�w��O<"	�?������;��5���j�/l�F[@�h�E�~�y����t�Nu��κ8���+� Z)C��<����nh��889z���-