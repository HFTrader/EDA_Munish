XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��G����_������u�E����y�/xװ�Ȳ��B��&4=�	
E�`U�D��`��>��nq��}�n�lZ[�q��L_�;�cB�y�o���+gM�_�U%s��j� $��n9�]��^�i�\��!V�b㏢w8�_G�.:�4�j��t<�蹇mП�i�i��B�� }�n�,7H�u��$�7*�P\*�l����0Y���=��.K,ű8]�oT`7F��]��>���z�~3���Y[Y.�*k�_N����ք�`�ceu?��Ț�
.5:{�O%�ã(��K�?�������-h�ܒ�����po��#��O�����T$�3�& �ؿ�9�Q��bB[�hǐ#3��,c89g��_3Q�Cd_΀Ԣv\ Xz���k�?:�V5!?�Ye�;v���t�ң]�[�bo���"���'���k����s�Q=�TU-�^�H����X�G\�����'p����K(����;�.?H��vӕ��>��*O��0�����|JepD��t��^fќ9���}���^p�~d��+�"<�k��S�]-
 �ϭ�q�prN�߹"К�p����f��G�$���Lm���d4�^^��eF*1��{�H,����Ӂx�E���L%(vd�������*��Z��k�U)�ϟjï��H��dg�y%���m�8��Y���?����K�|!^O)mR�ç?4�M�$@R�Q���l%��T��oI�\�4��;m�Ln�!���'G�DXlxVHYEB    9480    13f028	���P'~�]�����K������|�!�д��j[�_�t~D�O�E�={��B&�V��D�W�ւi���0�e+�~pG!�R�OEf<�lJ���6.%$u^�EA.\M��u��%��&�edq}9	t����p�M=�j���Sqfֺ�T�2�;�=!�f%/] EyM`3�v���*Z��^ c5Bk�O�e㈿��]�p��My4�4o>��O�eE1w����~����MyE$T`�$k���@���y��ųxM���D3r�;@<��B'jy��S��@��I!_X�^&�1[-��{z"��g��s,�k�Nѿ
z�ºp�oF�Y�����0�;�>�1�t�p}`�7B2O��d}�!���?K��p=�	�sc|f���T���u	����x�;
���Rd>��-��h�ht��$�tP!O�� %��Y�7��ޯ����`k*5�K�-����]���W\;�萉�|������Tȳr�{�����"�Q�IK��|�ʞ������Xk�蝃A��4WS��0T�1v�m��)"K��Z��Ԕ�O!�F����������������:�`.8��{�y'.�e���jM+ƌ�w�����n�^<*x]�'�/����Ɨ��{�t|M���I:�Z�m|���o��n|	�譣!�R�b��_W�?]$D��Y-c���&����R���;Vy�6�����s�\lt�+A�,�D���c�Ut%KcG�"iu\<L���A٦'��oВ�[E�l>��ܺ�B�2e�S��xbgᯯ�m�c�hv32��\�	�Oa���^tcQaI:�T����A׏P�ڋ��u-����栨c|���e�q��y|+�{�.�����:�bL��ض���J@�Ȼ���.e���#5�#��q��B��YSm|dyfC	��%?��J��b#�������%3ڠ���c>�r���/\�Ă�����@���20Q�@��:�� N�����4����*�[ B 43�,�e@��Oz�>��e�l0��Kوm�o(��@T'gO�اM�U��}`_L���LOow�Q�´,@*���~�op��؍>@�\p8�<Ƃ��_�VA����D|��?4u�15��n
�Bd��F�mh�OРҪ�J1/	g��3Ʒ�,�䂺�n(���7e5�}S*9[~����"�"b�5�>G�:�0�{�bu�\�[2����!�Fˋ69�Cb�W��q�ٴ��8��d(.-	�,,�0K�h�� ��s+�	�K�j�sƨ pt\��}c�|�k��Xp�G%|2�$����r	I�hKZ�?�T_�S�D�S@���TX�xfF��M>�`V�cZE��f�Z ��������Bo�u�9o��[���TO�k�[8���)�6��J�B��j�/<�L���H�sXE�)��)i���ܽ�Z�I>0ONm�ZD����Ép�ʖ4OwSiv��P7)��?`�Viz��K���_w��T�����(t�#
 xəZ�(� �1T��ǅ��U�K�]��H��sR��Pd"S����	��X�E`�=إ"���n��c�U�'y������%w�՗k��;=�eK����z畔��������1���]d�
�$UΝ)����4����L$�H�! d���`�PR[㹨� H��Ca!�rs`��o����D˶�������U۾���KFkz��6q�i(��SG�@ �������ϸ8��'o�91ްR2���Q���o�|D�J#�	�Ghd�]��^U~����?��A��ܧ���^��o�����W��45%�/�����W_����� �n��у�zJxxD�>��xix������ؼ7��a���H��� 6�����.�(��@�v	�ta��9>����i����*��e�r���o�}�����RS�-�5.���^^��Ȅ�S��Q��U�Hj���i�rf�ccKd1���DQ�ip�r�	��u�y��d���F��U],� �rS>
�O����fV;/��%j/�+q ��Υ�.`�����wG??�Iɀ[��銗 ��ty�ja�^�|�z�����FL.ͫ�4e��}w�@,���p&���u����Ԇ��d gy'~����L�t��K�Ȗ��(kB����/�{�D���2�Y{�6��
wʡq�b��DV�a����������ٲ#�w�c�%&�� =�	ۨT|��E�i��H�"6�hqk���[WăL�TA��v�`J�"��G�&�����$�cxϏ�@OA��v�ם~p�Z�����ˤ���Ў�Q�J6��7�� ,Y҇�}��$�B#Ʈ��/�|���|!a�9َ`���=e���б	�P�����!G�U�c����]�7�avG���9�+� &DF��b��*@�M%B.RQ�9���0MD�К���5 eZ����87huL��P��8t���V3�xq�A��xr'3�p���yD)�dҌ�5q��$�p����M�B����E�'���A7L�vKD����a���U��]���Y�	$&DO��������d�B�*.VD�*�{�-ٍ��Zz����-$}i٣�&�)�F}� �3c��ލ�k#�41s?��/Z�ӷ���,�6#xW2�s�:��RP)"���#0"�&��>�Io-F,O�2��13h��9:�"p&�{�CM�Ƒ]�+�d��LA�-��U��?h�� �#exz�|����0CKΒ��0*��$�W��R�{�+�d�"̊�D>���6=�#�<A����UB,T��[�� �qUs|�����7Ǡ�t� Ŷ�$@;�����_a�v6 AJ�L){�rģ!B�i�V*�B)���?K)3���gZ*2J)|d�%�A�5�Y�vf)�G���?�TUeZ�rZ��
aɔx4g �;禮��5�@ȼ[Cg�^����>D٦	��w�Ey���k�N�(��3�>����/���8�V
���{�q�9͉`���&>%`ٽ��~/+�ڷ�Y)K^S�7���$�*�)E��1oi?	��Z�1�%��g��q����^�H�.��#��OHvq?�_���}��V�"t �����<���~�Τ9rΞ=x4� 	����~�,Z:����״�ۚ����e���3�h�ܴ�^���eϏF��A�>�6��C��EM��f�����/D��=� �TE��NU��)Iq�l�O�«��Xe�#
�@�)�2�=���M8�5Y�i�������M*B[�����:YWĝw_8�e����H4;[�!3IRTo�ə��CF���:��Xڅ@lb���Q�u =�_���2-��$����l:.\����1�����	P18ɺ�k/��:�$�,nI��*dr���Gl�Pr�6�l[@��q��Ε|ԥ֓h��^9��u�R�c�)dx�����|Z�����RA�\Wи;��S�d_����v��4�[+UJZDB|�
>Q+t����(�B	�]f.�!��	'<fO�ב+ ���L�۩��W"�f���b�W�	Ԩ�0��ї�E{������k�������
<��T�/�F˖/s�܊��*��^��%�<ճM����f�����2󗭱R�<u������Y������������)�ܑ��*��	%	��ߝ�<�k�,�y�Ϡ���S0ѶX:`I�<�<�YGF#��vl����7��ݔUnv�s.���$8�}���;�C�-KT�\L����^��:8,އ4���Mg��$�s�s;6���F��퓦^�s,�v��RK�퇆!e#�'�=_|u�Et�Ҍ����*Yb$$H�~f:���	��p��5�'�W�����'n�aq�e��^�ˢ�>�������̓��[? �}���J���C��\�n��L�aƈ����7�8��?�t�����"�J�Cm�!X�c��h`e[y�.�Ƞ���M�S
8}��u�u��ZaB���s/��$��v^���.��#�icHf�#��F��e�p����o��6p���w�v�i�~>iL��	��.C4w�`��I'W���r��Z�H�F��U���X�W��tE��w�N�e��P|�,���[��8�򍆞	�)�n [�Ԋ2���㧄F��D�S-A�j{�ɄM�![�`�	�gxg&w~�T�y �M����>��\�B�ϸ)L��������V�����zN����ͪQ�%��~��㰯��4�\2V��� 0�j�s����@�����C�Vwn<ɋ��8\�'����yi����ux9���9)��,0�3�HZ�w1Tys2�Q�v��0/��ƨ;߾H�a���Ѧ SO4Z�-��O��LW�#_y����� Sn�V��7������ӟi`���iJ:v���<݆gP�wU�5�S!ЦS�rP��\��#�[�AtՍ��㡮�,�d�JvTL���h8�>iP����L�Ѓoh��2�z�ֺ��e�Z"DzS )U����/v�G��_A�.��0#��=�n��h Š)�2�[�f�A�q6�8	��aZ$�dƯT�s[����� 0_��)�[��1��懿=�������������;��?��ʲMr����d�` t
���d���c�z�=�� ��xoB�J�3[�N�'���O�h��%������;��y���\o��s@#��	�:�Z�i{bD�#�g��0��_��A�}��;r-�@���c�g�1�w��6����YX;?���V{��:�rв�Lu��~�����v9���!цz�*.�D'��y;lS)��Vly>�.��{W���ͼy����Yx���L�~0D�6Ƿ��
kQ�k�����JN4c dp��S�8>��:�/L���
tSb��r����MO�w��k�q����ͥ"mq4��.d�4�B�aF?�M�,Ok����쥶��+��U訂�{0�i5Hz��� u�Ta���i�<QU��H7�$PPH