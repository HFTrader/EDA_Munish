XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Y���?�4�x�#{R���8���b�
�`3�՞�z'�w�z��2n.&ۢ3��i)�t�+�t�	#7nZ���f�I��� ��p-# h��,���Lu#Z�a�l:S)�[���*��"V�!)��A!����_�-P�\�mFY���O*�h^�Zr�����W4�� r�^�!,;�E�#P97��B�J$���^�	7��)w��m;5�Q�h���ip�+���%����}Yi�|��C3bZ��}+�p�����lJ���>	-Q��i��u���Q�$�26��vPt�0����p	27����`Y�Y�5��,ܖ�u�%�`� R	���$wL�я%�ؠ�έ�!�'����85��Hm/]F��7������96���bS��@xTk�u|��4��Y�%O�@D�Ta}?�{�#��n�+�:;שm�ѯ��rbR����a�0��)kNH ���P+�J@����ld�N� ��P��!@�ڝ;�~;��%j�&�(�+Z�-K<�\g�(x��~�0RB�њL�}���!�²��<�/1fU�K�R����3���+��r~�qk�m��gg���r �.�Z�$k��Li��N�����M�_&X�1�W���mldY#U ��m���?� "G[7b:�9�Xl0n-8�;����Bڶ{Ѵ�r�}�2+�M�z>�/���`�C�v:�T�g$&��kZ��q������YO%	u�ѡ�˛���&Y��4ӆ �I�l!TƉ*)3S�ZXlxVHYEB    4a8c     ee0��ۢ�}aS��O:���,*�!��ܓ�ȶ��0�z��f�é�r���9���	�X��S�p�EN�|�ހcX���� �I{�(mv��QѨ�j�E+H�Z���q,�9�%'d(�/ic&�؂�;^�a�I��,��_M�kR��[b�>}b���l�gT��;
"L#��u�} {9�Tп�"!�ק�����ʕ�CQ�MJ�i��,
a�i�s.�¬+`U���B7�O�@-Qאs]�E�K�tr�}k�h*����4iZ+�U-��Id�ew0|V��� O�{Q�N$�f��>Yds���Զ���^�#�@�������]6F���߄��x��0��ɣ�H���tmvv)vЈ'�����ߖ�`T�#B��c��fO�袤�0sn����hh��!	D�@��d��kOR��'qx�o����yҀ>Dۏ&S��J5�( �b��W�dhm87%VNx�p�}~((���H�P#(�]�?�mjX�r��Y���m*�����l�
�m߮�ϔ���F>�C ��A��{�dT;���8�.���,3JR1`w��Q��F��}�Q��G�Љem�7�-�2��\�@H��ϒ�Y깨�7(N��t����%���N��1QP�]U��#��f�����+s#�FY4_E�H�l����]���~OQ9T"Ƨڌɳc����S��� ���Ǖ��t���Ɉ-	���C��1�"wK�F;��g�{Wv�y�'xҨfn�@�J:�R�^ٹՃ�2I�.��X��>�B��W�����+N8A�<ܲX�9�gPX�*���;j�ƶ>$߉?����;�W�_��&�݆��.�0�f�u����ҬQuK��B��[��CR�*�����p�TKyʦM1৿&�Y ������:Ÿ\�>X(@&L��*�qe�����]})	*�F~x�_
�#8tO~g)�G�&"���XUs�*|�w�jC�֌.��9�ڸ�3#Cƅ	�t_��;���0��:����dPiC����r��هPͶ��jP�3�s�Փ��6Vpp�����Nz�U�J�ʳ��q�$߈�y�A������$x70����8SLZ�Uw?�k�G�9Ҿ�Y���p\��2�'��u��Gt�I���Æ?��	�F8��cֵp�Z���;zyj�R?%��u+oa�b˟N&rdq�ܦϪQ<P���$'�ȴ�E�ؘ�]
����icw��|���3@ߙ9�/�O�d�\�D~�':�MI�ᔗ|��6��x\Aum����Т&x/o(���G�|�Ld��P*o\����i׫��5ٝ�Mj�:�!��r �4M�ʨ_s������!6��Ȅ8>eחZ��b|Hb�`l�e��n�9D��X�]`�&wz�s ��s���T�D^M�n��^��N$۰��� J�]�������mK�R±�{�+F:��R��`M�SU+x��ž�ǣOw�~FZ$($0n���G��Q9����?��6�	�nЖ~æ*�#g1�Ĭ_��&��NV��A��;�d�B��*U&�W�#n��EL�L���,!O�ZI#�S�~��H�)�������
P��J����;�E*���m=u[V�rh��}@�<8,@���3�Qv^r��R��z��h�2�vى�B���d�5�X��h��l|��� 3�P]ia-$������J��a��~ȫ�j[�j �lF�N��Kszڎ��n�4ux��Q^�,���s+s��9V��lNlլ*�����i&��@Mg�G(�������.h�9Q���qw�U/S������SS�&/P��	�F��z��εs/�kQ��2�2km�L2����7&���Q��Iꏻ���)��\pm3�#�R{�%�������z��7����$���������j��$I���8!!NW�7���$������)�$���N�MJ$��~c}O5!,��j�$���D��=�vݤ�f��⢕��i(�W����'+b��&'����N��6#@�A0Q>S��c��J��r����̷%B:����3��C�wsdV�Y�����m�a��Piw5qj�/C�t++1F9Ż�
��:�'fS�+�0�)�b����"�
v����;��^0�6!H�8;�T��\L��3M^h�Y�_���UA���fZ�5�n�+L�G^ɳ�uH�{��Z�9A]����m���7ݛ�9[;�pWE_�(�ar�Zi��ϋ��B}�'Q��2��F	\�rU�����趸�n����賽l˖M���c;�<�����bo�[�xU�jظ.Uz���5�}�1$͓@���*Q�'	�_t�Z�De� �[\�!�ώs�E�mF��iub�?����]�D���;bN��Uf	��M������\��dӺ��Z<'�6�dhK4��NԞ�����yk:ܼ���A���!�j@�+���"����P>�x6�F���Cb(J�s�W�?��
�+F6=��������^��C�+�X����+���r\%��1��+�q��a<����RU���ܷ�L����?N����-�D|pT�~2�������T���U�D,mn��������^!����/Cx���i�,i�b5��/GY��M�,$px!�}0d�c�� 0��\�H�W�#�r�#U� J���̳U���ɩ��v���oBD :�%o����'3tR�K�/�<o28�^'L�va@2�������@bXw!+�]b[�+2C�h���c��p����ݻf�2;܁��(�6R<��;H2*�n��'K�8�J݅�n���ƴ-���)�e=U�֗clA<(	��l���e̬Ik�D��=#��/�@���#�c�&Q^��^�4c$�Kć�JD�!Lr��C���kIo�T{��Y��#��-���k��|?�w�h�!S2h�/�1ˈ����
���e�ד����er�ӡ����Q��\A�ug�"/��A�Y�Y�Ƌ	x� ��I��4[f�D�x/F�Oӵj��hEi�s ,�N�L��x��|8�cF��G	f�Bz� zG9�b�;�Y%�S��{�3����	�Α�؜ոT&�ձ�s	`c��S�Y��x��v%�ȷ�۲������G�y�3��`���� �>���sC��$E�E��e)�v��vw0nC��"�y�R�T��@xNf�~`i�h�(�.\	Z�bs&u�S�Fh�!1Rl�% ��If1v�E3�Ԓ`q�s���(�df�Ϙp���){?�۫J�3�����_�t������V'i�;��Z֠0*|Վ>�-���v��{AXp�Y��9f|�.TW�����6�dq����g��nn	��G]=Ƿ�0����v����1���x.�&��8���#C�ڍ��_dԗ�i�BʴM�_8��k 茸-rIҠ������T���6�1�e�
����3��Jz��pKYվg�M|+
��<��m,�C�f�%��H�^f�{�-�F��k��x�d�!�r��k���`,.0�(#�mAp�%7��ꟾ��D!��)n#��Q`�<����}�T��w�B|� n*�-��y����B���T������d����y?�e��7?d����ͪCb1>�X
��ދ���#
�A��J�������U�,O�_7���UŘ	�v)�����^��E�x,�K�:)�C8��L���nR�Rň.&�6~�G}�ƂL�Gq����=��jW��>�Y}y�����J0��Comjp�� ��`���yc�i�