XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���j�8��?�D[���ГD�+'���|�&�� ��� ������0�zͰ_�k7����;O���iIO!yٶV�8{9�"Pf2��ľ{�4��+]������Vqq3�dh�D,��v�e����I}�|�`���M��+=He3�Krÿ��I�T�Ud�L }Peb�[!�Yv����+�Kq"s5&(�=H�?�ǌ��fp�y�J���� _l:��ʔ�����r�����A��{��qe���~9���H�[���B@<���ƣ�~�G*�0�����h6�1>������kRL��E`%����ww�ѻ�k�* �]����T��4E�@ٲ� �VДa��X*2�⢂	�O��L�jD�K.��~A�(�}�'v�S��{T-P�ow���ۈ�{zS��
{j'���G5҂��a`f*�5h�����Jh���{ӪG��HƼ9,�	�+������w���~S¥a�~�����}#e�E2r���j�D��h5���ș"-��<t�SEn�<��3��"�˼@�F�^�� zL����VO^�;3�'������\ �~�����F��$ڋ2��E`Uo�.�M��D�G ÞD\x|��?x�,���fT��������53!���5B���GO��Sm	/�՛�;A"h���k�+��y�|Z
�L���6�&��,��m:G�PE^G���}]d1�i
����ΆA��՞ۻ�|�hx��+F���v�n�[����"t9m)4��c�XlxVHYEB    fa00    1ca0�es��ˑ3swL�A.-���I^����95�y)Y�ULX�ۗ{Av�6s�-O>�OA�>2f���{4bF�"��C��������&�8���j[<\<�|�Q��LR�쏧nwJ�"��bʢۅz�7�����"��U]�(��:4j ��Ͳ�ױ�
h��n�`�lG۷]k?x:>Ko ���L���w d�����e$R�my�sL�V9$�n�s,x�5O��;:=�[��IKʦ�e����1/��o�������ט�%;������*-i]��"m	^d�h9#D,��S��H�f�)3"�h�N�G��2�'�@8:��M�4\μj����E��u��~��Ŭ.CB��mC�.;NחTµ��1�5ć���O��!u�k�Nhˁl��k�5�ӽ���
�I(�Hth}��=�_��!8d�ͦiF��ϙm ��1�e����]�+�t}�ţ���6xu<�gYFt�.��5�i	m��L&)P���z��+$#5��c��𾞋��
bkf������
ʲx(F[e ��x�7[�4�s�55��;��t��P*mÇ~ҍ3��[����U�UY����&Q� 1͹xσ�f\���x�>+q[���vj���^J��?rx6k��ٳ��(��z׬�G��X�.�����G�6 ��2�i ���Z3K�:,�*�e-`��&��=>�[���l���]�<��?�q������o)U@��:��ar�@t�c`��"w?+��F�D(O ��0c^	Ҏ=��<Z���vw�T���&?�}Uu�M:��;@�����1Щg�����]�����D,㾉�F�V��{HL��Z�"��/�έoTB���M�u]���
�YMv�}�����i�]����^�3_t�跒�5{Kd\u�/� )���ۡ��d=�׌��U�8�z�`8��n��lb�J��6��>eD�S֨P!��2�i��Jm~���$��ӄ&i4��+-���B1��[�U�T���1��i�Ѷ'��D~�ƭ��U'�cZ�s(�x�������N.��,���I*3��<}�����"����A����T�ܘ��Dހ�cDGVgߦ�Ƽ��A���D��
��\9���4�������mh�W/.�LD�y��qM<g�C�d�E듶������I�?���﵄z��oL6�����G���N�9�-iך�vk�j��2�_�|n0۽.��5OLd��hJ<̃���P���Hr]s5*�\Ր1��g�{u'���=�:Q�pj�n�I��j����#g��#�`�0��^;��@by���pq�6}x@2����5k���q,҇lnSӻb?�Rw�������c���jߓ~Qɬa��jXD���t���Ф������y��2jc]��ь�=�A!@}�0ӞR�
���`��{��v<Ӭ"�QCBTd�M&���xE�ЪS�!(�𦋄�@��E��s������������VAj��+a�yQ��ba[�R!���� =(eH��c����G.�-'c��̪P�����P�+���H+�|
]\�Q@�sK����]d��&�������e�B���b@��18���̇��B9�Z.m|�º��Z�X�`?OT����2����ߠ�-��QQ�w6����]�I�~9��&���Q���sj�eho���s!g����
��'������./Jj �\Bz9����ra�j�S���������X3JP���͒��	�NM����Z
��D�z�h~��%b���)�����v���*ZI���T�$�����8�5N����տ�Ƅ4���r��l֡}�h�m�s���5�
��4��>�e�m<��M�u��m���D�ѡ)����a54q�_������Y)�~M;��ZWa�k<e�R[%V����P�:�
��=��'y-�7�:}1'�K	(�|_���V;�2uj��v'�+-w���Y/>���CV�ۥ���r2����}�,���(*�wkVF�Sz���QԅQ�*׸����F�������H�]
a�����.nCӤx=h��M�ě��ٱ�}��}V\�,�5��+�d�ovC��6��PyL��n�3 pi���4��RI�P�1��|���e���#&7�*���w�3�D�ƴ���?r�"Y��k�'�]�p�2��>�8�!k���Wʲ�= �����󂔿K먐�Q�N7��	z���`��p�U�*��g��1���O��6o� s=2�'.�|U_,�3��F�\s��`�E#|���#r$���ڨ0�9~�LOF��_"����ƈem	s�!3�+Z.Q��K
l<��%$��B�Ca+����z�q�l�j@��2����b�U"^ٞ;5�}��ړ�Ϗw9�Z_��MQ��<ɣu�������Վ���e�Ǟ �����$��ߜ�,0p��+ࣗ��>���æ��{��6�\0x�H��������)�����w�Iw�����W>3&�z�T	ܙa>�wBp
vN3i��D�y�)}�>c�]�}���:�>�����Ux��S�Ю�!�y�̆Uby�~�Z3K~�}^�U�].`<8�I�I���N����'@�mZ%{i�,4z�� ���C�S�pI�V�鈾"���!���	2;r�8��h��_�4��D�꼓�>O68~�����+y�L�N�'��u9W�ҒxK����y��~e�5�vy=�-�'mo��������&��C�Ӂ_�8��� 1�`�/�����~�}|^��^�M�eM�5�@�M.C�"��s��VE�	M�o�Ə��<�4�`H���-�~܅��4t����:�}
r[$��V4R��[�����S�DFC\�7�`� ���oHA��	c�7t��_�'�&��kKTOތ�.��R:�Q2��F�BE��_
�vѤ��>gֿ�=y�B�U5��	g��6�"��Hg�~9uLѦ=-`�O^g�o%ef��@r٪��3Ds�aG9������I���>���UŹ�0��
ȶ*b����?���.���_Xt-�'�y7�N ���q`5�<x����L��勺��c:-(�k��W*z�~�{|�:��%=2��X5���.�}�ÜY@/��6���$�&Z�0���Z�"�b���;\6��I�>�a�>p�-�\�d9:�`�$�L!9��Ϭ�t��4�!3�!��zMc�5^�Dd��5GT�..W������� �8	�cib�:���<Th�n�^+;#�5!��؂*�@3�y��H0��gF�s�Ún¾�5κ���~�4)�,�2��d��5���A���`*`���ma��2��¹k��Q���o.�3f��ػ��)�@M���n}|�hP�a���;zX�B�m��2��Z�\1�#���mu�s^�ǔ�0��!�GIV��mۖ�{!������>���1-%�6ibֻ�=�m[��Z��4ϫ�;f��'v�m��/�[�j�!�0?�s��xi÷�!���<3�4�	R�\H�_��>���+ �����a�Wyg�Ĭz_�5��Z�����N �wk�2jf��mM���ȹ�}-�.	���#��&�i���dG�l�eS�~f�k����ЬӦ���A�v�
��mDb'�YS�T�:�+!��4�z:�*w�wX�w�0�y������n!p�O�2�&��"eX��o���1BV��Θ����^+��C7] �D������@$SA�5�x2�/��|�}��G4뻘k�q����[EP�����7y�)Os�l+nҋ;Q>y��v���z�8���*Kl���2GN����&�+8�K��	`��"�PZ�e�	�;�`��P�O.�P��Rbxu"a���G/�T9�(��}���Y��vxs�J�t��tx�~��)��~���웏��nm�4�R��dyC@;Fq���ݛ�ϭ9`��!���� S5�H���,��	�7�$��K��<����M�����/ٽR+dO��c�N���{��M���*ן^)׆���V�8,C���q��eH���m���>.��O���[S<sF%K6dX�=Y6��{ d.�������X�O�<��h�3� �4g ������Ziwˇm�«�V�?u�ó{�eAI�3`�m�g;S�#�*'d_jR&��x���o��p�F0{^�VLيVh���$����7��m}q����K8���B�7����,^ݵ>!�a!����訷8[�io�I�^!�L����gP;*q�%��i��J�Ó؅���t��O�Mp�R_	�ao$��9.�{G`~_��5�pәM٬9�wV��2�75C%�$�X�d�%�˩U>%�yf�n��5��f1S^d��o���mbsO��?ϐ[H�Bw)%l�6b.��֟y-�wI#�&�2��R�,�b<��s��������=�o݀��4���fwG�<%:i3�6w�cO�Йh;�� #�X`,4s#R�י��d^�����!�ބ+���@P�.`w癿%fEO���F�+������3+�_�q����"�s�6
��ɐ��s���?��1H�	��q˄5� �׳���"�Co��
�%��3-),&�Nv���Zg���+mZ�54d��!+;�9c�˂5�,��Yk9�حd~�W��@+B���оh�4g���B�y���K���_�>�7�TpF~@6��泓uO�~ţ+����S����3#\o�M�����3���Bp���O�+aLE�vIu�M�Z<�� �սNqhUe~?���E�>�����[�N��0{��ﯝ�n�][LW�4�%<u�>7��0��進�O��Z^�9�Bnaq�R2^��b���k5��n`Ӣ�N\J���\�`����6����<�Ȯ�{�긦�dQ��tH�˿9�n��GaH�������-�����I:�bq��쪼��.�
��!s�r�1��Xh7�����_')#��'p�Ɍ���묳(�!�(�t�����p%����#�3'��f
���^^����Ry��Ǭ'l��@⸑6������a�i3E��1��֦ؕ4*"ϥ�:L�S
��E©	��`�u
����� ��L^����Y7�I�ܬ�9(�f������'ҹ�]]��a� +�w'��~9O���|�?��ok�"���Y�J�;��}����BǄ����WeI ���3�@��+�}0���+7�1�6󕁢�U� A S��ۀ��4/=�N9�S������Ʒd�	�}��Ki���ȏ��b7��h�搣�fv�%�5za�Y��y���^�Q�a(�r��c����m�4�/��U�<�� �e�ڕ��Y�k�!����-��d�Hb���d1"�����%!�O�/x�-\��W��9 H�����#�@�6��ag�L�e�܆�����ݒ-�p~ƕV��J��KŪF�*�=�q��ԧ�Q���S�	o#�/�����Ơ���K�x&���6��ѻsj�(kP��: ��)*������6`���B��t��;f �|Z��*��/c^��ʨ�}�9i 3hLH8����f�Gf���fhd���b��|Fp�MB|�.�V��f!���돦9'�m��ǖx��0�f
����3���*jP���5022�iRp�gL�E	�xo����@u�ٖ��?�?)�=����f%-�%��'�� >�[�]�g�m������b#WIjU�s�)��կ���.4���=�-�jǩ�d��ig���#�-
�
���#<~ʋO���P%h���brOi�}���@�L���^�3��|=d���I��H�:�ҥд�nyG�I}7���α�a��:'��B��̱=7���-#�Eؔ�ɩ;@����m3Krfv�4W���9x��ܗ]7����'��;�������7��nK�x��x�/���	��ܓf�£ �M��ͱ4]�[�� }`D֖
�]�c�5K���
�8!�BQw�d ��E/��}��y�c+$�0��%��s�T�l������C�gU�E,T�n (��G�c�k��A�#�����Z��<@��i�)��m���m��y���ω���[nU%�Ա cyꀣ�݀��	9<0�a�7K��\�U���W�iN���`-ֿM�V���S�H�i���#^g����0\Hd��R���	�f��uB�
��`Eq1Q_a6��heY��$cE��/�8U�4)�ibZ�z0��%�@/�Z�����
	,ܮ<t��J�{Y�4'8��k �8�f�OG+{�E8�r���}�N�.߽���6Y��I�Ѓ$��2|�M����9���OkZ�kT0�����k���2"�q����PP*Ko��>3ԓb�����kO�J�+�cۑB}�O���m����@��|k�hC��^!
�T�P۾��ǌ���-c��U0O6�~�#��n�N7�a|	_`��'���kM�'��^6#A�u<a�ϳ;8Ӿ�w��$@��ƃ;� z�R��QϚX������g8��?���.Q��b!���u�ͣ����j����[fh5������C�5e2g����K�th�foτ�����(�`��W{��V�0Y�G��*W7[ˀi-���(k�?Kq1�u}P'�uFs}�V��&#�^�l<��G@���yJ�s�~�$��X5�E [AY]2���`�d��%��]��`��g�-�Y��o����ߙ/��t��\s��e��	(t��,a&�~��J�0'Ύ�:��6R��%�ҧv�c�3�mS�U���0������F���qYBB���,(������<��hܒ�=6�ܝ�]Ya<���M\�2ܓ�y��o�j%k�$���}����9}��~)*/�.���g!�,��4�Z,.S��)t�Գ�D��<	#o�	Q)8f��|u[[�cSku�`9 ��W��啸;1q���.ѷgT�80��M��np���R/QI�d�$�C�;
 Z9�H�!�ӗZ�5����	Eטx���c�O�8�_CY��7j4��]&��y+�BmB�9�T�A�E��U%
E4qX4�y����j��}[�͝�O5ͼ�~,g�d%3�ZI��n>�;"��x��CT ?4���tf5f_>Пg|�gow�D�x���c�w��ܞ/�� �*L�-k� ��X��?,�uXlxVHYEB    fa00     cf0�.��c�ԵR$�#N��67!�Y�%�����D)= ޙ{J|ty�͉sԇ�,+�ǎ+T*��5���B����{lt�����ˇD/Y�/y)@��On�Kv�w�Q,��w1���:�G:��{�@wl�n`_�³��m�h���:Q��1Gj����;�-���49!&�@�u$nb团(F�j��v�w��ep0|�����OI�%�J	�>sb��jx��Ĕ�JV��L��2U�S��ͨl����$V��2�6��*� EJ�p�+4���<�I�Ƣ�?��<�4��1.�;/�Gw���l&��6���D�UA`���;�~�i��=��m|�w�.r��e�ob�=�q�D�_J^zl_�ڨ@
�.P�ޭOd�9��+D�#�] E�v�LRH-{W8H} )�aZ�u�J�}�~���ܳ�j�y��]㙕�Vh
Pt�l��;�(:�59oD��e��"��.�9�_���T�}Z�b]Fn��`.~m��1�
p�0+F��*�}�����.~"�Z�2y����ZT�������Tl	{���Zɍ]-�����x@" �����_" eا��LK8H)����_n't��� ���s�u^���6�g��)�Te0�t~[���&����h��S'3��'40 ������J���?G��9��O��8����G&��=��������L��i^���/�)��U%����>�8���ŠD7��I
�wpc���O��TH�pZ��4����NC�A�o���-�7cV���s����%�*6�QX��?>�H+Z�3�q�S�k�I���w�lyz�=�ipemx^,p(�]|g���C��;����xG
Z"P}�/����	 ;�Ȝ:"��]���s�� XD�O�8kҺ��ь_�K_Ϊb��1BR����z�}>ZZrR5���4�����)=�I�@%��g�T�4�����\�Ф���f(SD��y�L���4��!�vЋ��i�U�i#�]6�d��l׉�Q���Z�ւRe�%�I�h�����#�="�����0�W�ӱ� ��)-����	��r�C�/��X��A�|Q4ɣ5&|ע��{�q\Q����C�,桜(�
�&��l�����-Z�����l��=`
Vf�ǉo�����z��z�Õ[��`�{I��=����,���2��((�R���i�2��3��.�~��EH�;D�J���B�"Ƣ���c�R"NeuٻdDv$*��U��tU�O��\ل���_Hk�\޹Fc4']���B��2���
#m��@��˼&!O`WF�����Ģ�������D�;!|n�I<�5�v�c����o����k����{߀b�vc���G��<���&�b��Kv����5@rY��/�{�6���ôn��� �ʀ��Q|GP�L+��˛�P�w������LAځ�pqM�*��w^�!�@Kî�*�n"h�k�N�u��-|AZ��B���{����	���g\B�	�'o 40��t��W���;�PE2�#.I��2Wғ�H��� ѩv,W�q�%�Ym+T��O�c�^��gtw>$�F�����\kp�#]a��e_�[����Db��Xq�Oa��p�J�TY���d]����d�0j0ܿx�~�ݮ��R�G��/pq���1�l����xl�H�a�B&��&/mG0���(��������<�"���S.Ռ.z�TS������խ8Sn<RR���������T���T�����B�>A��{�,iZ%v"p����}���q���r�OV&��A�q��3\��v��|�Z���@��@'1����+DA�$&
S�/���X!7����V	%[A,�3qJ?:���c�,Η=�U5�\c)y��p{�(gY��6��'���;�L=��iv��Bk2>
J;�U#��8d������4�˟�S]�� ���:��WtUX��A�������8�,3�P��叞N��?�z\��D�HЖ��IH��9C5����#��5�`0��y�GSǙ[q�6 8뒤��[��/�T^Q�m��d^^�ϥi���ӻ�n�L�n�O�0���J�aW�A��N�yV��Q�X�x���͈f�Is�)�m���q�"�滰�7�bM��\��ԕ�٨��-�oP�5���ä鉄��D���	����5������qA���͹���G�I�	����!Tb�C�g���=i�D�?��@]��nZ��(Y^H^�t��t�1�}��� �-"r2i�\2#�A�s\q���(����������k����ʣ@�C%%��G/y��tB�۽	�M1�K�I	7������Q,1�C=�z���.P-�P7� >f�ē�'Ȳc(N�S�X��C����IKN�
����b���&B�K���C*�����������a݌
Qc/i�V���� �W����"��X�	�s�=���O� Gآ�}*C�ں�I#P�ª28������E}�⓱�Y��� dl�>��z������{؏�G���5R���y�pR�K]��l�|U���D̆�T8 T��S�刨G��<zWu:�q6�G^L�DB&�V.��>��	x�Gw��&B Y�t�{�[�X��X�̹iq�;͸��"=!N,y<�� ���C�,���"�G}J�qJ�v���QȐ��$!��Ê4������ݴ���c��X1�a�U� �f	�(����v��"�<��*��L�un��c�Uق���v_z�K>.�h���<�����XU��H�����B�}�`��������fa��Iх�	��A��Y-�� Űt�K��:J𡠺߾��E�*|8F�Q
vլ,�C#���^ܓ����%6��6�������P�j���SUV���|������Ga��ϻ�b;U)#u��ZPl�F{|`&����*\�:�k�w��F SrR��̳��c�����9z�����x)���N�!gM��#k�M�"����jSI�IY�aw�2d<�M��+v��F��Y�0s��tdZ�⊮;'GvΝ �������
�m[�l�����w����A��O'��0Ӆ��!��{/�q�$o��r�t�c��Ψ��4� z�H�K#�xǕ	N�!H�3D�6$:Y��<���yw;a�s>�6$6�G�nP�×�Ɨ����sPP���a�C�4��1<�%�(Y������Wc�N5��lC��(���ݹ_C	[�;f���6WYf���wa�1m
踝6>��.�K���%) f���^n֟XlxVHYEB    3981     4d0���Rp� eo�eX�/�D�� {��j��,��^���	>�B5��F��_���R*�����;`���鰛g����Z]7�!ku*�� ��9�Θ7W��_�^��s�3eh�j�ˆ�%���*?F��[�6������
b;x/zaS��߃���|�ɆY���z��[|�J?&�'a3e��r��T*�Kל���yڇ�aȏ̟��ٔ<��0�ls�9�xƵȳ��L�sc�.uYem�E�%1� �������h=����O�����/�~�t���'\H@k|ad'�r�!Xl�������z����짶��[���+���U��h��,C��s��l�L|H��Q�
AV�5�b9M��r��@Ik6��VN�-�0-�5e�Q����C���j��ֈz�毭D/7T}{3����6;*R��-(����Z�m�Z"0��ɭF$�J�.�P#�@��p���u_�En���t���i	�0�&ۂ��Z�8-^� D��E|��h��ɉ�.:�*��+�ӌ6a����۬��V��gE�T��l@L���<h���tԮVK�O���yӫ�D�)�X��D�\G;����ふ�e�s�݈��,�
�fwWIj���9�~��)%��N6�])]��"�s�ß��D��W(z5^��-mM#A�?<���H_�V7�6	�M��'/C�l�|�U���բ�{�[����i�3�w3[97 ���fN ��.d�D&�TC�u�﬷�PV��ʑ�@�s��C��wd�����Q����Ɖ�%|��K�����2wF�P��E���%k�4cm.��b�P�E�.rG�kZ5P�jh9_Nt�-`���}�k4�ZS����U�/yo�nV�f��-��iQ"�ǐ���:��M�U4*�̡PN�0@�V��hsF f����zcX?�j$i��W�F��?���z%��aZp���"�ǳ�����ה���?����6�гX��=�
�������~���V��>�F�,���%��j5z�cA�J��ۚB}9�;9�t@�_����`�����d�^wƓ�t�����]H�/9��
���B��hZ#���W�'5a�GCF����F@L~&]RDP>�NJZM��(��.�g����_�i����n��3H��J�8���*��*�o�Z�*�RY�ܧCA�fvv6JXP� N(��