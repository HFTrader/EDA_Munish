XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E��d^p6sX<�)nu@P�i|�Z1�ƾie=�QYT��aF�8�baz����˺v+f�І�F��.y����	��A�*$,��B��5S�$}��yj#�y�Ѓ��r`����W�;��~�?U� �?��y1���[l�J���ܡ�����O����4O�AZȐ5���~m�Lh��{I�[�F#�����������j���@�汑�$����
/�@��e_��3=v���D�i�pl����Yk.���~1>s��_�F&B2S���5ǀ
�H�ߨH���1 A��N���Y��")�[M7!HN�[�K����f�����0��idP���2����$s\�r�k�.}i~im�vɨ�/�Fo�[� h�h�^�jI�	�7��D�qi1�E�g���e�y&�~52��R�5W���7������!u�a�jo�V��r���kJ�;�4��;��a@��E����&S?��6zyIl-�@�c�l45/�ȁA��RK`F��v�՝B����϶��gc2i�a��f��B���i�Wb�x��#�.%��I�)�n�X8��@�o�	��7;@��981]{<h�EM�mg�A�1�����o
.o�SY�U�}Ȍ=�ۧQHi�n|j;� S�[ޱ6W9�ͻ�ISb��;9_qAiӌnz�x�Z���ÓG�qI�8�s��a��0*۟g��|
��/��N��q޷:�����Պ� Ryg"���j��ve��XlxVHYEB    fa00    2040vw;0Z���a�R�.r#r7��Eտ����߄��枞�K�/�,���V����ޔ{N3�̩���N�'�����ێ-Y���3�#�]iW��5
��K�ub�g6�:Ef���,���#y	=���#�0�.U������>��,��㓈 5ࠈXW��%+Eg�a
�}��o���)-GՑ�tI�^�EV���v�e�z�w�q�Q/���:��M���"_�<���K���s�.��/+Ð��F�ڜ�)1�X�ZK���K~��3��{P�:3&�ԗ��>v��Q�Ŏb�����u�@fYO�8��D2��d�=��{>�)��ek'=����+R�JL]'����-B����1�t��	eا�%�DD����IG�
�!޾4-�������,K�~����,+8s|�1�[�DPdٚ�Yv+���{��+�.B�҆m�M�Y�#���[���+���QcR�|}6k;%����XfUtZqeV]��Ƣ���Ƃc� 03J�b�~�E�WoC%�zR |j���ǾZ�rA��m��d���<]@/oe<����R��#?�F-쫲�X���R�\t|C�P0�E[�y̆������ �s����=�XW�1%�q����:��ͦ�m��4�l�??�g���W��m%8N�K@��b��މ�[�etI' �i f�Dw^m��7	�ѽU���+hw3��̝7D?[�q)0I�,�,^�UT%N���\P��H������N��컃�{����_��O�v��x@@˩iA�t{�sP�-��KC��R���nx��	@������Sj����s�@��Ұ2�UUǶ�5D���>�L�"L�c����T��_OשŅ^5����/ŤR�!ʵ,?�+�c�~��aW���|�A���ne%1��E�C�x����7��d�.:=M@y��7�9in��D\6��}tn��e��SF������$����L8� ݔ�B���ʞ�4&���c�F��7 �a陷�yq3,�P#~ ���q&qOf���l�.����af0:<��������]<�tۺ�㶒cb�Օ/;�˜�t�D��Q�1Nm��`ZǓHpT��d>	�% %�>�+>L��7l�ڃ�$kt���#t�@����_wd)A�4*R� J���2��6�X����D쒱�n� �E��G�w{�1� zC}i���j��
�g��c��>G���{`���1q�����l����^}8T{Y꜋
�P/������~�s�׌DH�MTD����� ���i�4qX����������v@� Y���N>�]N��"�f��4sb$`wS��D�͓��+��������(65�K��&$Ϲ�u6�"@�%��]W�+�.�E���ˋ����[��	M��>�O�[��{+�k	�}U�_4�JP��&��K�V)��+&�N?S.�q�^�$j�ͅH�_w��h!�e &q����r`8�c����pX��"H&A�{^��$���M���{����z�6�~�����z�n}%����8�?�*W$'�#F�5T��D\R,'���G�𣟓��b��O��R�c����h�� !1�%��w�U�YJ�u������	��iC@��
|��.��2챿�A.Cj�J���������Y��`��0=䩬����
2>�ѧ��T�i���>ֈq����9I���庲i�x����e��,�hE��ɘ6�����졷���ry<��p��۴�[�UF8�Qѡ����<���!;�s5��������Y��K��-[R��-���}yQ�Ae&�@f.>��;=�_n����X��6Nq
٧�Hiby�Ԥ�Gr�R���ç�-���赟�d��H����)��m��vg]{���ad�(n�ڱ[O����/���k�j�i�&��!K��Q~��:#+%�7�A��QiD�v�lj޵�tZ<�� R���%�Gk��'��D��*1�X�s`�y��0V��+�7$³��'oY)��|�s��X`�7?k��vp4����dS�L`D��"�}[u0��|kG=L��K��Z<�.���y%n�Y[���>5�����G�r�gG�	�z,�8�od]��4m�{2��3�X�Ti�Ʃ�m���1ϗ"��/�A]�VI��:HwE)�!K�"R�KaѾ����
�|l�O��,	����L� �?���b�#3��׉z����8��S4Z++Ľ�E�<�`j]
;�濦L�]h[{@��%��sed���젵:�5�³&u'�h� �؇��R��+�"���N�N|�`�+�'�����SF�u�2���^i�$�^�MGV��"?R	�Y���h�
�����9����������x��L� �p�}tD�֏�AwͧRS�˦O�J�P�g�Ñ귪��©�/���X�A^Tw)vTg<r����~�sF�!�����Wr�z&�.�{�U�TҴ6��;Qa���:�]Aw0�Y��m�|�w*�C���?}|��擤/1�SD��|����+���w�{f�@���jin�I�4ꙶ��&��"X���.�I�hV{�+d�����(�w�w�D:����	���;�� *	��{5rn-�H��[���:����c�.�s#1����	�I�k���I���=J�![��OD��Y껙ch.�>8�Rʈa���NH.}�{~�0{$ Tf���74�7L:Q^x5��IR&�0%�@8��-2�v��L-�x�Y+yL�'�@M��L=�7�,y��J�
��d��om(s	�먯+�r����f�q�b�_��8�]�`?��@��"��1���҉��:I�M���HX���I��0��*�����Ɩ�1`%��G단�a���S�G	V�w/����{�et�n~��,q�H�~e�����sT�O%Ũ����U�&BW>\�u�VӪ���~��~CiA�A���[�!��&�+�r�}]FpC�a�Q3b ���9�`�u�w��28��]2�{�i,Y�]NèJytT��ic�	���⑃���4��T���N�
p����N�XGp�Q�Ϡ@�q���-<LS�����1�5�����'$������T��r�	�y݉ł�2*l]��x��\'=(���#)�:C`��82��3�l$s�)q��ɬÙA��q�=������APPT=�d�p}&��;ғ8�XR�q�#	-}u���=�{���BԂ���n-����
���m?����+:-�'A����2��l�[��y�H>pr��7r��j�Q�F�נ^��ņRf 3*~�B' ���v�����Y�xø�5IՔ[��*aST�ҜB�j��P{��yV�:<A����l�G0X6(Q��+y�+�2����m��szu�n���ڇ+NW>_��D�?�F᥍n�J#�&��ޛ9���V��l< ��dܡ�����}�|U?M���@�A|���w#9�^��P;L1�x(j���O�vC�6�I*3f�"�8:p�o�u�rP�h��������Wm�w�";�7��J�Y��c��L}�9*da6���W�y�i�n֐�	Q8����T{/G_���4���� �x1C������gLΉM�p<áL�Q�Ũ����KB��x23N�k��ボ��)�4�����{Z���R���@���|2ۜ*����饿z�a��b�괔R
\�寮Ty�!ӇT����mD���<Yr�]��s3�^d�-X�-�+a!�}��Li����������l�=���'�Ʋ�Z��%��=
>�k�9�|}�X́�����o��6Կ��ܟ�D��ɀ=Ȭ�k�E9�rǋ�NA{ð����8�X��m�Dp0����O��|��f%��~t���́�c|2���-ԴC/��*�{|���=��#�0O7n��Ƥ�BX2\�c���mь���
��@�c���u�2�H����������s��������'�ũN��L��iCG�Q��1����4�xr�r�w���d�Iw�*?�=N^�XZ��L2��/��2K�%��f���0��Y�V=�0����ضa^�)��#a�T@���{��J��� =xCҸ_��\Fz���2�p�)�Thg-Z)V6�k��-���nFr���|�ޚ�y�R"�0Xd����h<���HC��HS��%�[_�G�eY"v���L�M.��̡ݸ�	XP�S��?8�80h���ހw �h�è:~_��Fؗ�Kr*�����d�j���c,Ƙě.�rYք��Ҧ*��>9��T��N; 	��=���"6AXn��E�L�D��0 @\�������/�+��n��u���L��f�za��v�`�=K�)�c�t$����S�!��Q]M�Y�.��\��6ImyjI�|s�)$ۭ��DU���횈��n��V�q�Y����KC�`�q���xa�(�lFd'�f`�kvC�s��q�u�k��G��\�������D�~+!�����y�ZR��J���:�,>�7�KK}���<�^�_��y���n��W�α�~G�y
�t�ؼn3�'e����6�B�'^zBs�3w���<Nᙉ֐��բ��Ua_��C�~�X|�+��zqNf.ыeBoc}��J�~U����wi�cY eq����ѵ$��g��TZ����d��]�S�G�x�M8�R#wy{S7�_�S8;�AH����~bSt���.Q��*�wh@�R��_�G(�.�G�j���8���v��K_ {��"���B�7��s&hup�Vk�7�2M�����t�3r�')���5 �����W�{{�!� �Pi���K�����m��_,�VU�.�����d_{lA�V��*X���}RK��i��JH�	��`Q�~���O��8���ԣ�ȂO��[��w���be��tt��Qܤ֘��
��*��5ȏ+��h�"s��{:����F@ ү��4k�S��wf����J5-|8���x�ip�աfڈ�O=V�y�?���_ط��4�C U�H/s�)��f���We9т:�w##G�VB{S�c���]�� �ɢ��(�@�B�k�����9(���8��1���chj�W��<\��Q��Ң��!~��0s����HO��3L�[ȗ�-= s4-V���e��2ba۠��D���E��<F{g�ިڄ5��z%�m�9P	h�4�,?��5�����;��NPL����WCN����לz����i����G�6� ^��jpE��N�֐Zw٬�A��H���*����O,nj5�X��s	�3O�1y��.�����N�V�H����Ór����!�6Ӑ���6M<a�LޠX��MdI�(,��W#�_��r�����5���x���wy������C�Z�o�j������@x�|%��-3ؤ�XoM�/��u�
�)�|�l�2u��0��R�L���]T�G�Zi����~�.�5:y?d_�)��7�0�VM�Rב ��u6�Q������9�$��?�;�#h�	2�,�-�/C�A(J��ęƋ�F!4�TS�8o��"�@��9�c�6��K�vF�]ʔ��ؓ3��/��+s:�t=ڪqNtΊ�^��d���D�9��CHO��8�i|�^���o51�se�m��w�.΋���w�}ׁ�y�|i� uڄ۩��o�s$>^��+�+�*����w�p��:���=�R�����*npQ�PџB���w㴞h�h��x4Hҙ�D���\��a�@Ţ��j��o<G������ǟ��&�E�z� 0�UY��(* L�So��?%"ڶդ��%<l�]����� ���=��z���ڧ�N���k��ѽ�!7{��nB���<d��&���}��%t�]<�b؜���E�W��G�.�AM*"v���
��A*�1� ��B�7��{B�)S��z�܆d����.D�z�ÌC�F)�G��F���1����K�+�g�^S���d�L�Ɔug��j*��̪x3��f��#k''�C�Sݟ�*Tm�Wf�ܞߔiÀdNF�(^:�}�zv�I��qcv`��!�Y��C0I_�x��U�2��d/������n��م.UĐ��τ�~��*���4���d�1ҋ=��KC���6�j &��Q�~J��Q�/�wJ��WGoӓ{{��m �b5��]-"��G�4�Zn�Ex��	���������Z_sxp\ƴ��6�a�u�%~� ����3D�I\U�D���ۯ5�&'�*���*3N�:4��<̓>��,%{�?��*�ԑ�2�@��Φ�,+N�8��f3�_�Rk	��Y�Z}t�~5�D�����c\�[�T��M�v��y4��Ԑ���$36h�ݩ���ş����Bi�{*8:�T�����?���71hL4�VVe;o��'���%��˹��}2�Fķ�Y/j=*�J𵰑"��]͚�+(���n
����7�[�$Q�@�]$#�ɺ����5:��Uq��*�Bk��R�x�a���ݎBّF�!�=sM�I����\����,yMHk4mG���مz��I9ϰ>�=��)�󘻂t�H٩VXG�Ҫ+zk�TG�4{�B9������y�k���xk�"3u�k�e�Y�6��ch�t�0����;K+*X�3�%�A��1�B2/͝��z\��3F�w+ExM����s�����°T�4D��̅�a�늽z�_��`�^a�SX�!,���Ě�y	�	l.�$K��I5A��9�o��f�9�tl��]�.Dc�R��l�BΩll	�U	�)�Q&���Q|�u�1�2���QƯJ��A����n������]ư �!��p���y�,��3��{�_9� �d��)��mݼr��|��� q]����>��;��C�j�HKk�mc�Q����Z�لrվ����d�X�{�[Eрa�)����1�N�)����:�,O		��ۥbV,IdY���(���k�T�����4˛.��G���7�冭YM��ez܏����pʒw6⸜@@�e�Rh�?ry譾0��4����x�)c�O�i�
��G�NMg9>�3��rÃ�wgU$1i��B�z�{�[@@����ָ�Q��"Y����$�J�^?>$�� ǘjި�
!���͘Z9�u�Jg��.ly�I��n������O��I����v��o��67��^�A
6��B���_Od��$x�����Q�y��σ���5�E���d�$p��rɀ�Ϟ�MF��?�^��6G^�V���]y�j7%ǈ���(��h�wm���>]я�b�Z+�y��%��!�$f�i�L���ry]�_��{@�>��*J�+A��W��p�?JEu�Ǒ�0{�9aI��F�[r�##����1�tr�G�(����J�ެ��kl��'e�R�H	��%P1DL礭�Z����U'�{H��v���k{s��� ����fT���;'|t��$1>v=�M���&��x�����.��;s���!)���)�i`�1�ݭO�R�o�S;I�������cZ~�O<���u�l� �b	��&���9ȧ�ٰ�%P�!�H����>�#H#�7�X����pz��/[ɞt�9��Xu�!+y�X�u����RQ�W��@�C�h�
�p򤊾�77עv�e�w�D���L��=���6u�f�3���2�|e'�"��i���cw�L7��h��9��o��A�l�2{,�|hb�i��<��1��o���-v~�`�e>)U�Qo0��Ľ��6C��(��9�aSpH�0o�95U���8҇E�NнҬﴤ�E<
.+�^"Rq�}w��%�a�$YK���݂=���g�R�i�0���~5���x.q>	Ga`Z� N?�U>�K����?��rB1������%����A���k��S��L��m��t6u�V��y�_0~�zf�p�[|�P��.�6k��&w��l�V�[��;jA��oN})��\����H{�:���EN���<\(�N�Z�=tM�4s����S�Q_����SJ��.�@g�UTֆ�S�^J����ߞp�7p�oV���*�*=v��*�@t&���yFXlxVHYEB    4f62     b50�a��&�s��R׎Ib�(3g���2�E�Sl�z&vu�k���sY���Z���1��<�퇓��7"��s�n&�nmG3Q$3b����xR��[�]~�!�8 ����g����e�"�i%��ݲ�y�GSay�}U�(cJe9��u0��V��b�'.>%��s�iʩ����0�n=.J���Q�!{ds"*��\�=&���B1�,���:���K��t�����^b�R��7U3�޹x2^�U"�Q��,&[F��ΰ6���`Ln�'�.0W�v�.W�JQHNP�o��6c0#�]#�hz��¢��V�/�[8�Zh�Oc�x��c�vy�+as�����=��;ǡ�I~H�l��D���������ʍ��@����N���D?c�njⳮ��?���4&վ��
<PD�ʔ@����+�o�O`ʳ��9,���?����	�Ugbd/�N���ei!����������mWeu���ݸt���=7��T}�a�Q��� �w �Z�2Oӓ���_�6��Ro�������ں��u��l�Rƀ�G�{ϐ"������㿳|����{�I=&�a���hw�߾�:�_�-`�9�s(G�/!������^�v�3�?��6U8�u��U#�&Ͽ�js�pڿ)�����à�1{�ي�e2��a۱�2U���#�Y4��3�/��iW:B�/z�|W8i3:��X`��أ�ffp��3�2^��@����*�	�k�xca6��gG���I0ڗ��
�-����s9M��E�G�/���DL5_��"�7�!��~��L����[�5@��̲6?���譌B�t��+�d8�w��X4q���R���>��B`��?��hű|�2���i�yL���IiKǦ�MN�K�qx���m�bۮT!	��C!	9���%X��k�7r���uu��#ۡ�u�����4�p}A���$ҢƧ^�� 5�<����/M��Xn'�hN�#�-Ω��n����0����2����L��%���,2G���"��kntw@�z���u;~�c[��=!Q���|��MY�O���L�7]�p���Ǳ�l@L���ٕ�ljI���۳�U���m�z�t������Q�Ir�x��j����Y-zd�w�6'���5��Z�U����(��ʝn��"ţ�Ee�&o�iO�n۔vț���Xh��DX|x���%x��;��w�.�&�c[�.��wV"o��iS��O���xR���4u%���h�JB۩��s�vI�-�?G��Z}����@ \0�O�o�C_-��GH;I��>��OW}�;G+CZ8�U�!-h��O��f8+�2)0lo�����iFQ��"�*rk	dI%F}I�ߟ��@�9�o<���g3�lqc���ঃ���냦��\؟2�z����N
��߰��HH�P���[.=]�)����H�J���TP�L-�������0ۚ��s5�E���ʠS��5����
q����*8)D޸������:Β�=�j5����S��,��ǥp&���������~��7λZM�G�����*�\>V��%t�AZ|8�������ۦ�]�$�߳"ml�E�}�{���j��%VB�=���dJ�oEM��m���.�s�yR�C�<������ i �*�3��	�H���z�Y5h�3'%��T��+�Xu8�����s4����X_=�+����J�$�/�3�ǎ����6�w��+^��%�ű��x��D�{6G�V�}�䐐�nj�3���q������킬zfF���0��نb}��(�qf%�v� �<r����VW��@�X��}͙��h_Z��n�!U�`�uwS��1|u�Y4� ��8��d�M��ws@g1�@;Apʔ������[uD�t����ޢ�Y�}?��X�}�e-ٴetl�s��g�$��(���(Կ=��찲��"4p�*�.��>"�O��Se�]K���nI���T��Է�������Dfc�N5��";d?���a���+��?e�qrԜ��{]Ov*�]���C�K� :gC��k�V�nl��Κ��NJ�EL	��l���\�]�E7z �!�\{,�����󘍑YJ9q�iԂ�-4�B(���~��k����JP����ڸ_��χ�.�~ǖ�� ~j��4����؞�1'�U̩����[u;�=�I���w��@oWs�5��f�¿�`���#r���-GIϝ�B�����_�
��)�O*�&{ ��A�2��
Nm{Tԧ�7=����	�0�"ݱj�ѡ��ܺ�n�&���B(�(#H�\ɜ��޾1�d@/>]Ad�9�/��H1�u�QL"���p���+�9!ߵn��{ٞ�'�{KDӲXY���0`{�""�$�g���7�d���4��Ƶ����bp^����Ҥ�Vc��(��%�ܞ�!ެ{�4�z�g�L>t�a��#��l�b��s�V�~���36�)ky�}xa}#�BI!�=����R���5}.rvLb�ϝ��	JJ�A�5�#�x���R98�~&��Z�t2�XT�1|ٙ�K�����w�������u(�2"X�P��h��X+��Ezۙ�����I,�HVt�BIl�-g��r[���7Ɋ��%C-�(�O0��$�]��ܘ"��tKwh(6_Eg�f˟nOE��nB���:����Ҹ��Y�wG9�������%�u��u�>����&ڀjX����a\��_]I��O�i�#�Ҳ5��`�jZQ�����v�����k��v�R�������@�b	4]������/�V�|s���C	i��QAyQ�i�Z�{�l�9'x$��c�