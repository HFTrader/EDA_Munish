XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v��<�l���I���C?y��f��J7����	�m�]V�Q�u���G8�Y8���2jn��ϓ�e�4I�)�92����{�¸1=� �YoU6:���79𸃓�&Ot�n�p���
`�7�}�A-.���1W���K|�qĠ:ĉ��2�|�*��ݱ)5�Ӏ��*v��[j�v`�o�S�Ty�Ocz��6��\���/���k����D?���'(���<�G�����e@��|zL~	4�e���>�ǅ�ЛW��{ �f�Fn<8�yNaGQ��!��pAf�O||_e:|�w��Y6���\�M!�Is���;)����$���zm�4ʼrߢ��me�z_&�9?�qօ�Z�˜�6�x�ϠͲ�S�=�iգ����3� �"�-`�1���4���-e���������ZD�zK��4D�(-Ey'c�~g&U��a�@Iy���m'����X���T�QI��K�<�����mb�>�t�����'�����16��O(ڱ��|��MM���mR�ww>���-W��r6��ؾ?�\���뱪+?9�_vr���@yJ3VO�Lұ ����b��t�E��|�z�숃�j7,���/H��>Y<����,n��?�3*4����:�i?j���r��`�Y'�)q�"���j�je{�^e/���qFR��i^���=��e��mNDV/{g�bHDoӏ.�=��/�T��0���T��fkC?@�=[cݴ�j�H�f^�����漢��$�XlxVHYEB    5df6    1510Q���&h`�n9:��T|3x�H�;1a�O.mp}���J2H�y� �AJ�+�Y	�W�N�
ln�pD&᱋`��i�����^�k��n��P&���W̨-_�w����(�%���J�_C�@-3Լ�`��B�q�-�
�y��:�Ԫ��?1��b}��ZJ"��wm��:5�w-�U���#�1{���>(!�;�S�{W�Y���g�B�H*�-���6t-��<`8М��/&L�����N�PhQ�0��|�����Z��P]ܧ��nZ<7V_�:��妿ƿ�(���I�W?�gѤ!3�����
�� ��c����sO��=��(�6:A���G Pu2�Z�|g���sY�������Yf%�f��lQ����3��DڔFKL1�����@��N'/I�x��Pu���n|&qn�s:�q�Ys�q����O�o�š��6������z
83qZpX�:��3��I��e�m[?t�m��}��I��c���2ﯭ6^��zD��]qrg=���d�o�x_] ��wy����*W�.u��u[m����������>���8S�A*�L�贠&%E�q1��0t�%���E>�G .�1��h/e7A7��K��-�,d��sq&	�����T�6R�V���)�l�포\g���2\[L�#qN&��1U�Ճ�ߦ�j,MdK���r(���,�d2��;2c�>��h�2gE�׆DL���� ��M��9�33a'����K����w�G	�k[��^%ʆz��?I��j,�-|�4j#��a���\��Dh��n�u�8�h��V������c�|4���#V���������,���'�Y�D�tKQ��I�j�v$#˿�
l���-O����\&#ӻ�^w����ܯaE�ߓ#I�t����fQ��#_�8!Q!���^R����pa�J�0����~wd�g)O��ȴ���Ҍ�-�v����S�|��D&�uD��$�;�q��0��8o�NeN.\.; Z���W��t��m�3�'��{K�*1F����JG7Z�T�㨒Z)���w�;�m<�F��3ҥ��^Ðt9�%Y,R���g@�E������Ȝ
�M��
'��SG�xտb.�z\��n���x٣���
NpA3�2�M��LF�I2�gj'�[�ćM��6!� Ȱ�e�,�CŒaf��j����[�%�Ʊ������-�Ω�mATMH�~�ᶮ�`�֍^�;�Lw�sɺ��N��{W����g���蕮Ökc��=����f�wg"����W/3�V�98a���BOI�8r s|���Z�m@�����@������3�����<�S[�D�;Ì�ӝ!{X
�G�m@Eb�/�D��j�����4}��Ē�"��9k����%�?!?䂶�����5Ó�+��j���d)�;j*�-P ��ʄ
+
9H�r|���l�����HO7�(�N�KM�zƼN���k���a�kL�r���d'�w���t�zQ3�D@�/V���}A���A�J�qj�NXE��v5J%�"�����N\s��2�*��{�]�B[$k�:�䘪���RRKY<RA5X6�'��Փ��К_|� �4�*�6�<1ڨ8�5fI��i V�����|O�v˞b������y���H-Nӿ�?8)t�f��	���nh�γ&uwB���V`����\7���nB��R؎)sݭ����c)�縅��F�����C��s .a�0��t�8��M�lAQ>j��/������CER�SL׍��a�K����i	�a(p�ƌk��X��iU���??��z7��N�'�2S��Nl�L�T���ST�9��+���gX�4�����F��R�[�òMH
*Kw����0�w���l���r�L!zR�vϳ�w�^�,��6b�����h
���PV��OC)��={���x��� iH�7����G})�����ku���D���-��^:�q�L��������Ds� �ڬ/�9Or���8�*��O�IC>���@0���H�[�Isp-�f���C�m��Eh�`ݒ#-�~���F"���uϐ3P��ӈϭ�S$�Z~������������A�#�I8���p?���-���qT�C�)�t
�
b�؍�)4p�:h�{��I��>������1�g]�l�'@�	�˼x�l`�M���Ð��)��1��tDZ�8����%���Sğ�����s���L��h7y����Q���}��(����%��E���9R,��Un)��5��$��aa#qL���+�XĠtr���8f������L��?���	���FT|�_V��[I�X���"�[�-�����T�5���'>��׹�>����V"L�/�b����	�D9(�A�р�<����;LM�����x��#��	9=�.�S7���v��1{�6�҈�K�-�M1�����Pɏz�v�����YF�8��J��h�G��/�B?�HnrH
��hNO(-�|�YZUzy������g8�*��*��2�"MJ�|�6���؛�4(%�����TmɅ\���	��Xv�^��R6�ɑ�m�����t�^ u�����6�(��[
�-���q�r��6����=&�O���暻�������$�Zj��e1������X�.��h_֥C��A��~I˛ڲ�׼I�')��D���a�{/�f��9��W1���H�bd�����ZB�9�l��bR!>ŘO������`���VB�|=��g�0�Ǎw�=��$�����+�|��1&�@�n+W9o��@�`��'ǡb�c��jK~>��}����@s�9^�Ӧ�"/�[��&j*�rq���Q޹�ܪ"��F9�-F�4�F���	�Y�$\�Ϋf�g�nWLo��[�ګ9�����}�Q��*�->��jP�9S�-�����k�s�f�CG���s{s~l-^N��3=^EV� �3�O�9SN9 ���S�4�d�K{Z�?E����8 ߐu��?1r���Q�k�#��/��͞����L�lr)0�Q��i�[u&0�����B��G4�0K�=G>0 ��P�0�w�3��#��ᓩUVD����0�|���v�xdg���WLꩪ=X�+ט��� F�9@�Jgt��_�U�u�z�ۭu���/�[����iDys�^��9��7`�,����{*����pT_�����a�!4�ͱ0�ٲʌy?�I��� �.I�:h���.�� �.�\����}���k�)<���4S��WH����6ŧ�V13�LpB�7;���o��GH�;�a*e]O���g7���PJa|�r����"�G0���͒�t2j����X|IN��=37z]�)v��yk�^6��yI�~W��JC��*�eTj�` ���9bGࢳ٧ڌ����}UKTR���n56)Ȩ1���6��k�`�%�V���VA�)0L�YHm�b�o5��#B�}�V���J
)K|/�7is�DxS�X�F.e���e�>���I�¼Mn�+�e�ݽ��RR��W����Z�e�^���Zo�E$��m�oj\�*!��e�80)L�X�I>����娈)~��I36]Q���"�B�~�+�$xj�1-�����6@��O���}@�����.]��{��̿�7�D��n���2��]���_73� [�8s��]yU<�ek�x-y!㸂��&d���T�9�<��f��1�k���إ�(��d��%ЀGQ�dKS�@���)�ǿ�C��:�|��V��u��G����2��:)3Y�:Y��A����f!F����o׽��Yd��pf����zdٺ����wĀ��w�ٳU�FG	\\>�De��xi����,<�8�6 �&��w3To��Io�G�o�����cx~��٩.^Z�n�9w��w�H�������7��޽s�.�AU[�@Rm�[^tRm����ƿ��0FVhͤ��e�����ّ=@E�{�f��}�]�C�� 6�w��E��'>�N��!�D%��b�g��ʨ�^0�9)����[0�el�FHth	�0RS�)dql0g���sb��WFNux'�@���\	0�.��ݠ~]{�ƨ ��]j �j�k#Ռ�k��h5P��и���(�� ���Ua�ύٯ�*��ߒ=F�M�&i^�xw������f@�@�y�E}��5�j�v�C��}�7)�B[��5U�6����0]=�aK����9���{�ǃ�n��ģ]x��>2���$�6�Wv�&�.q��s�Wx�-�����]��:���kWFƝ�ߛ��b{��I�{]?��������v�*�b�[hԒmH�?��Q�p�--���6�`���%��^���<�	��+�)f�3�L�z�r�c���kI~���A[H��G��5ѥ���	��gm��h���G�)s}���Fs�k轆4�7�p�вm	 �1���^���k')E'=��4�3� !�B.����;C��/�T��^�����Ɠ|W��%�]5������Rc�:L��/}�e{hK�Zݥ'w�5k,���3|+�@&[J�e�APY���<=�F���/�ԯ�BvaI�(�<��]H�,̺)q���w�"���SHz��7|!T3y�Q���5 D�v�E���U�&7�J�V`1�eN��)~Cv� ��l[�^|B����jA+j]]�
Éw�d�%�7�X�%CC�5J:}�~����������Ag�
��{~s�����E8X�H�x��������
Z�* �
[V9�)d[��~���A�0��őj8i^X̐H������<D��d�6t'ޗ�=+�&�c]��U�-o
�L�T�Nv����op��6-��~��t�5���"^���i������QF�J/@��i�]�t
X�N�@�o�i#kz��#c|�.YPL���~�ěI�
��17|��p���.���<����}rmu88�^�{��F���g�m�(U�a��td&J�T�a����ȴUs���|��SJ,��O�V��E��GkGO��0�gh���,�����7]���r��lG[�=(��7�&Hw�y�]��"5��i�ŷ�q��u���x�i{�{��sx�G�����%���+74�H�w��%u%�ӌ�����%?g�jT[��IS���h
�F��a�� �Ҷ�G��4B�ш�(e�w9*���-�$�(���+��7��$�A׋&����z�؏-�y=�@|0���D���eC��T���9l|��%���"ܦ32��}~�b�-P$��	�e���ٰ��d���