XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���o��z��(�D�j��W'~��'�ƲB5�&;I�h���ri�����_C<	���&�j�2��&C��W�Ga�wL��n��"���k��T�m�e��0O�a�ខ_��V��v�>�jP�@�d7��tc�퍪S���)E���|�����`�i�F���}��O�!��Hk��z
�Ԓ�~��5���uo��Mk�3K��m�(R�.K�!r���[��K�V��e��05��,:�����@ն�Mf�;?%���\�n:�8#�c�I?䔹�MeԦ{:��N��Q�?0p��HJD��ނ5���Mf��=�Ef���':��Ĥ릅�&m�I�mQd��Cg�O�>�K$�]�5�ŝT��e!Ćl���jE�1���HHG��G��j�Ι�G-
�-�����yO0XLvg4���z���(�HD�i�s�&��g?,��ե8����N�ʷ�ayW��v&zG+\�C�@�0��F����[/�u��yV���OX��+i>4�҇��OH]]`-��(�����I�4�#Wf�� ��ⷦ=���&ҏ_�а�R?�ZE
��+��������N+	�>.���*1{!2׎�z�]��OB�@q���!�B�[�� }�f���(�T1^�_6XD�(9s�;��x�'I��ЧgC -p�gDN�L��ϷC��z�;�a̾:1��2� �,�hZ�M^,yn����㔨��8��@f�4��)��fW�Ы����n�7�DV��/�}TV�wXlxVHYEB    20a9     a60K��03��AJc�ɇ.)X�-33n���i�����d������S���J��G����b�[��@��ٔ����D t4'��2R�*�m�C����b%H�K�2��\F/�@��@�`Onx���D����&�)����/N]�/��^ a��8��9�v��8�8ؘ�ٌ-���ƒ'Z
W�|-I�/�$��}�:+�,�C��ޜ�E��X&x%��s�Q��,�'$�!{�II�
��o�0���a���N����l\��^h��sk�m8��Xg��-[*{����5�_� |�G��Fz�bgZ�H\˝aY��2�t��|�� ���$��p������*����G�_�A*1��e��if	*%���*i-j�`R:������J�e>���b��s�q�����(�����*�T&ؗ��Z��?� 1����b�L������"ĝ'�TDSjb$�������Zݤꙮ��[n����P�ݜ�*�E����M��X�!!��|
L^����a[�gFS�$6��.|�G%��.�����	���m��#��@u�0�2f�$y�Q�|@w\;z2��Ugp쭘Z��L����7To�=�ڒ�(��e�4�l>��`�B��Om	��8��X.�d�W��$[
F	�ݟ�s�DcZ�rɑၬ����0�J��q |XhJќ�bп$�_V&G(hf\f)�<�c�b�8��:$I`�:���_w9s�0� I��0�W�_�0��:�˽b��ѷ#��L`�{��V��K4�i���@��^Tw���� 0����"��e�5%z��e
�9���&g<�?����O�gnTЄY�Rk�p\�2t5�d���ϝ�B<��]�Mv��L�;��0��9S�Q��a������T��,�i+,u$�p�jޛDS~�r<�:Ōo;����	�=F��	���������1��0�p#ZmXWl��S�/��#����F�H����U�rģe_dr�2���^ ��mE��M���I.v��6k	��ܐ���/��3��UN��u�(V�IoS>��Dژ.u�[��*t@F�Wd�6ɣ�J��N2�mn�f��	yr��ǉ�q���(�������,a�!q�4�����@���,ш9z;Y�Q��2Ӧdϵ�V��4��狢�R�%�w�"X.�<�]�z���>��wD*��2�9p��OW�4p᭤��R�lT�o`x|�2Q�$��\o���)�.��:j^�L�_Ƥrެ��_�t���C�o!�!��ZQ0��	�`�/.Gz�9l��+b�R��`Ҥ�����y(�̆4�B�^S"G��Po�T���g��H<`+g�VB�Q-Uwh_F?���S֢���Ja��:o�hS��_��p�ɐbb�J=b��Z�SN���9�D:�}��L��V�i:�* _�����H@�	l��N[���F���n�����9�	��b�D#�O��	��1��T�?���{ˑhb^����F��`N�U�D;��iT�u{�D�ʠ�����:j�!VC�C������%�=ΎgcH-=6�s�n������UL)Oeʒ9�
f�Z�)B��@�������Z)���Z�x��G�V�'���m0v��`�_�;v{�,D��󞤜��eK��ːA��߅��;~�I,j;����X��X�+>����3��LJ������έdT�*��]j�?�&%;B�.�ƅC���o�c����R��n+ �4�q����J����僖j�("h0��<��(�g�	�0XR����X'��t!e��l��__��u*/P�4�k?��lkgA~tS؎5�6?3Æ+�p��݈KFci �).N�Ro��|i''xB9�)��Pq,ǎ^:�M��N��^gJ��iR�I{�U�ռ�ӧq�{�^��g��2cb�� �Z���o�~�
� m�E>���+�g�����h��T� �-���}f��ʇŊP�82��Sݞ:z�a�(�i�s�Fw3��XW�z�[�6%A)��7>�ًxѺ+�Aa�E���M�����At1b%K�6�I������i�g���"�� G�||��<��{�8�m ��a�}�JE זJ!WX��h�d�$�
�t[)v���1����oW�b��bH�O�w�7���"{�����8���AU=��y,G{Z�@��MH��`��zH�__3;��0�ӝ&��O����U����0Z6gD	��0)_�,k�v������;^Ng�::�rd1����,f�L��8A|@�7n����I��Ӥ �Ȣ�
x����z5�k�%�{Hϕ@u��yS��^�?-�vݧ��b�Exc�7��>B��C��>0�s}y5�ЎQ��>����T���~sr��������$gK�Q;T�R!;5V�^r��W��ba�}ܬ�NJ��|�"�A�+� 2��h�?HRŖ���:Tp�hi-y3�vj�B�����/�ߏ���of�=$k�5m	.���L&.'R��a�*d�b�`<¿b��� @�7�����+0�����{�����r{��>7lѸ#8��k��V��i͂�KV
�ǋ�c������xX�
I�ݝ�$äD!.�v�f*���iT#vB�