XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��\5��i�X��Z)�B3��"�(#���`gK��J(�-��������*�0�� �芽S�t�o/��'\vd�q.��o�?_�<�ጒ��H�����9���XIb����D���k�L���G��f��gm�M�j���Q�(%z�KW Z5��mm׆J�͌g��߲Pu�����n��~A�����uH�RIOկA���� ����vKVj@���Q,�p.�b$�-�Ӗ������hby�Tx�<��d�c�9�q���i��,fX���_�K���P
ωL+ǰuƪu O�� ���|Z���l����,r/�`\�+�f�/"3�-��]N��r3L�.��!?}�#��)RK$XvKK�P��ѫ�>��,����x��Ο,�>%j"�߫���'=��+_�-��R�AWk�=M�����6$���Y͇�3�$|�8��ARDc�z�������\�c*x%@2�r�����?'�QH���:�����z���1��7�Wc~M^��Z_i�FGo�$t��'HJ+�_��}���q�+-|��J��6���<�d�O����U�� �c�M󽊫FP��ls�Dc�D�~���F`��Ŋ:��.v3�ӏ�a����T`H��d�?�)cfG1�'y�ך�WF�T��Eٍ-�����Hn^4�-|2X��1^���_�#���������͕�Yz�'������o�u\9uD��G7�h�����ʮ	�h��'Q�e�,ȥ����XlxVHYEB    1da6     930�!��4F����Y�Ako�;?�t��Qfv��$�\�^�䁀�3ӟ�:�C�<�H������@<��b���W��o9�#�TD��&�+�{ն\�����WA*O��Ia$U�/��Æߌ�v�A�=ʀL����~́|�3�����y�� ���C� ,Ib�į.�1�B>�}�Z`�R<]���\�ޛ9ʧ��f��������2��}s�¿�;MǞ�-�]#������*�d;ி'�<@t؛�±�<���MI?���S5�����wp]v�
�E���l��R���;���M�\��K
	*. {%�P�Φ��l����I�Ix��̲�޲i���Fԥ�[� ӡ�j��o>w��`S��mn`X�&��ڸ�?`s�I�t_�*�K�W��.ُ�����]ٮ��}{.B�7%��Y�n��^��&i/4�ټg�`"�V�E��[��n��~��V�V��GL�ns��p��=����=�K*�?�
����-��v@�#�3�2<E����(����"XҐU�����-�׹܇��H���Qc�9����!(j����T�NVj��:�;ic���C��c�EЙ��^,~z�I�ɵ��be͸mj��C��d����T��p�?zk�w�Q���A��d���`�qASu���u�p�-E??�d��1���+�҇O�`ՇS���a~���!�H��7���]�I��|�R҂��:҉�'w�o:G��y;
"�*�l P�Fq�m;�c�!���q�f.[G��޸���-����t�%p;�iL�����m�p�aG{r���0v�]WЁ�O��3���)rRo��a��Bt����lz�����\���λ���ß�S�}Y{�}X���Ȅ��o䛱��'��@#l���[�{�+���é);���(��ei4��0��$Y�UF	6k���%7��9U��9�Zb�i�|�|����*|�
c@shPQy rU�{p={	���RN�D�;:�����7���̙���g�'T �jo�-�!-^���"gp�ö��#]�iZ��[FG�1xq��.��?�8 ���M&ϸf�N @�Q�~���j�Qv���Tq��ᑻ�g�;m7�4_W��>�6&TWnX��Bj������}�������8��疗�޵��k�9�e�{~`������nm�7��z�^M73��Mf=_|c༓E��YF��Ѷ���yz�yA֎����󖺀�^�PmzJ�g~Fa����
�WD1����^��	1� �[o��!)e����J�W��Ѥ�k�Zȃ�;�<9�i��P�B�?�.7�~�:��:�M�(]=m���f�'
���B&۔�P~�?���,��vLG��F�3�ۡNR�|t��[-�De������t�K�q_�����v��h9�v���o���������!%��/���7K�i7��	~B@�,y��!n6X���Yi���ҋ�Ѐ��j�f�β�J������"�H���y5��	���9k�(x�֟����ߗp�!C #�'b0�W�x��o;D���=�>Uk�߶*y�<J���\y��z<.G��B��N�B�AH�G�[@�-���WC%ds��{�Gȏ����:��c�-<�L�dmu�&��q��T�rԃ��`�^�Z�c_�+��<"GW����/��É>v���61����v'��Hz�s��l���5 ��q�CB�A����h�'���6�j�X&�P+
�W�Y	��n;}����b#�LR���E���p��f�ىˊ�a7ap�z�_�"c�F����)�ח7>�*��@����&�+Y��4%���%m~޿ߘⲞ+���of�[����m��>c��4����0!���YE5�	�K�"`��Q�qŖnM_�9˽ŋ��\��C���aO֓kԆ
8����0oZ��q��A��p��,��P�}�k�����zt��_��V�CB�20Yr��K�.��$�,�{f�,��?�#q��������l�>����o;����Ds�d2��ƍ���$C�Ѳ��8�T{�ʠc8|�������7�%���SW[���ю��Et�����-�QI(��[�݈P-���M�9��uǧv�b�w�vI���XwP��÷a�
0���z�s<z	�dD���FJ"/�al4B�u��@���1n<��4Đ���_��׮rJ�Ͽ�P�.8ճ�=�5� '�)��8]1���t}�w$����ڨ-4�kU��u��c����솥E`*��v�mm�e�%2t�����r