XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���5z#5m�c���	I���bC��p.?\��C��m�"��a� �}�j��;r+l�	#�a��Ld��Y�_ƙ��oI��-9�Br��i����4BYVYV'��]�,�s�w!J S�؋�9�5v��ۃ��ٵ*�ƻ��U��^�!g!%9���XP���(;Se�b��+Ç�@���B����*tΛ.��q���7,���ٷM��\"���+�N�+��7d�"oPOsC���0�k@\���ǼW�%-�Ue�'���$C|ꁑ���q���^�W�=�r�����%c�z�RG̳� "�������Ybn�1��0~Șz��ze����ux�`Æ�$�D��c�<u:�H��KB���~ۅ���s>��f��%�L67�.�h���zh�ZO�"�Z��a��[�\�޾;��^z��B �n���k��:��ե`Z#�(z�ǅ0��x�Vmyi�.�cpAfx���4x���h��_���_[��9��@>���w���Nqd.?���)�u�6�5T��Wz{W���h�C+�i��*�|:;���yœ��6�cp˄�B�2�F�@-�?"A�77 AO��'h4u|{e��oX�+ H�x�r
�F��Mg��׋$��	9�QX�u\kG�l��vT��|a���gj�Ё��ꗆ9,�h?
q}j��P�V3MK�T��D�Uf@ݼ@��d	�8�l{�hB��,�[�v~�(d���'�O����P���U�q�\����LT�_a�XlxVHYEB    aa52    13d0q_�t��1lƯ��ݿ��@�Ǌ��]�󪡙4�Դ�%�_��WǸ�=�!�ޠ{O^�Q�ǶF �v�v�=��ݭz^�kPǆ)zҦF��c������1Ց	��e&t�i��WA>�-	�Ҽ�*p�����_��H��9�l�(����O��YK�Yt-�p�V��I�2l��wXmz���8V����u��ZY����x�K��(����/�����ӗr����p�F��;j��P����X{�U��+E��%������+��Ε���Ç�����(��#lY���C�V�|���3�BSfaD�� -]]�r�М^Oګ|��0"tj�)��V�R���ɳ�@8@~�}X+lyK�B�|��������{�`B���|��?l��4�w<Qq�66���7J�8��-!���*�u}P�lr�M�S��?{�-�Y�7:�pT2�f�b��F��3{N�?�0�L��CR~K`Si�pDN��@Ma��;J:��g/2}�z�ʪ=|@�|�py�`�F��Bt%��:1�*v]{"��sXX�â�A�#5� �#鬴�E��ܦQm��(Xm�o�*ˣYI0Cwk#�����	� �S�S�vj��g贊�⨒�s:���;���š�������ǉJZ��9�}��Φ�C��ŕ��D���gB8I,��x� Ȓ3GZ`7,�1��Y7�ϒ97�!&�h�;��y�KW�:2�q�,,Vf"Q�������! � ~�ڔ��.1�=�Y�×�S��+�4�xgRԀ�B�ca
�S�#��pV�>�tK��W��O39�R�~qpJQ��7ڦ���j#�j	Y��Sy;�J;#s�M��GϭS��zf�>�,�����⧶�X�:��������i6���AS4�~���K�o�x���f���e
�.��+v���v3�^i��uO_��8��^B�c�Sg��dBg��$�:;���9�ud�?H���JE]i׾�����Lo��Gr*��oLg��AS�B�5��M���9��}�BY�QS��l�ڞ���"XO�g�����<E�+�^���s��w�{��Y[�گ-ԃ���R�]uT�M+`8Y׆*�X��Y�1f��~�ʟG���,�;r?�
,�i!J����)���7�kBc�PG�P��8aB/���ڶ��/N�*��}æژ����YgTPJZ�p���I��a�y�c%T�(��`y���O=���۵sC����Ü�ON���+�q|G�AXX��v ��Lm��T����av��s�Ѣ����e3Wzm^�Z |�fZ"tp��!��ڬt4���ץ�zC-�!Vd&��IL�P���?��Q�y�������R�wS�S���/|G�)b"�2p�^�^�mR�4� Z�B���uw����K��A=)�}Ň~���~Bg0��F��b�c鳾�%UWk^S���@MWQ�[�f����ma����&ӲƓ>�k�L�v��(����^�U���Mgͬ9�5��gYl�E~|���I�
��-�O��G�<�M|1�`	�}����
�袑=ɹ�����9Fn&����� <`�?��������p�c�����°�~N����F�x��05cXz`����V"|�W���F6Ψ����S{�c�4W��oӦN�ODq�fI~�)���zn�E���{���N?(?�'b�I�=���[!s��J����H��L�(�U���ǣmsP��h�T#�gG��/uM�Q��&3N��"��2�G��X���3�=�+��iW�?^��z�{�$׵$)�*"w6�u���-�����r�D��Ky ���>��DL�K~�t]F�2�m�Խ�a�U�</�o�J?�y�����3�� ����u�`�=�J<k����f:oZGI�B�>:2��F3*U�WjN��W�����І�~DHG���Im.�N��e3J�)���4q��(c���GTC�
Uq ��{ ��w�G�(��C6�h���S�
�  
Cp��t�I����rH*��G`���q�v�zBf���z��\���r;2�}r����! ȉ���+E/�m�� -��7ާ�� T���\;B	���o��G���v�7)��844<%O�)u� ]rD�8�,�E�G��u �H %Uh������4��������6��<G�m�e�`b�d�������~�H�����`�����M�2N^��P#�L(�A�"�s�q����`���Ox:�t���F(�U-j�:~�x�� $S#��tU�r����	S��6zg�>ol�#�O�ZܔʛN"&'�q<��8��q������'������AGC��0�}~���⩢-=�����SI�\��{���m8
��B����ѷ�FTeZ�[�VZ�XL��j9Y�T	>�9h�u�*.�
#��N�k�)!�#�̋Ay�����U��ȅ:ar�j�'��@��tv/x�5b��Dy�&iOq�S|�?����X�,��rE�y��>�9�i�B��҈�]����j�W�5��~�^9L�DZX;�*�<�`��J1�V����y���,jX��Yӣ���3i����e6x� نb(7����ܵ
A��=X�k�����d�x����VU�$6ϟ�78U�O�-]o
C�G�z���ts=S[auX[�bs-���ǐw�Rh���[���|���Zd��f�;a�;)�W�uډ�&d���A��o>�0'"V\H�6D�e�Z~&��T^�Y����@1<C���\�� �"J���у��cY�*�A?3J��v@v^'� ��ZZ�������,	R瑈�O��N&l_�W?5�6����Z��M��O�B=�,�іc��	�`���Zq7���E��P���ֵ�{�0o����C�Y��>�@p�s�R�m'Z���3BNR�����،���(z�}�;���u�~�_~�h�)t�����چ�q����J�&�=��/3T~�K�<��˗@�,�6��W�a|�f�O_D��[x��j.�d� )�Y�Z�`��_8��Ҍr�-���l
]1I0��m����KRnv�x��҅ЯU�P�K�����(3;��EG��>�E�����H�E���@3)�,r����t̽�fE3�w�C�w,>����w�@�e�����&��;�EF_B�F!�fTz@o[3@�%�㹰e��<���M2�R۔��U2���W��"���$��"��ݛ��:�CK�]�ȹ�����~q�{�׵�U2>�A��'�7�Fٶ���5�f�����fF@��{�E�H�e�i��Ԍ��ᇗ1�j�aj́� ��-V�a� ����<ω��Y��߉g�6\�9�t$�/��k��<�==ZM��N��Aj����Ԩ~Q-f�d�A��,�P��~�'!�(�H��L`��Ě�B��Y��>dN�_N��6_��5_,Ʈ�FJv.�K�C�K��(���8e�C����]��Q�}Fbqvb�	�_˗I?���4��" %& %� ��M��FC����O�u;{=Da���R���$<D�Yz �o��zV��p����@�����R`�ݼ�'վ��A��C�ᕇ�3¯?-x��l����Q.�C.^�	g�o��9�� ����Q�N��������D��H� ��
�*'���I��,d�I�I:E�w�|�ltf{Il�بU�$�#ɹu>�/mꨉj�Y�J"=��D₄H�&C/�
�CSp1@N&��<� s��%6O�eK��Fa�����
y�R47����ٶh�zū�����5��iN���UG�]bn1����+v�+7d`�	.etp*M(����%	��ttj�?Q���]:���M(�5U7 o�o��
7��>+��"��A|Z4��
n�&:�|+��>e�X|�-�i���3ڪ�<��
|����+��i��y�$��(!?�3y����Xu���d����J#�u�s�ٟ"JX�u��~��SS���/�R>ɵ!<v�-��pJGNIa��k�)��WA_/i��*��kh��X��'�����92*,��%'��N�SjR�Gt\Ү���$�����+l���et;������U�BNX�@��B`��`s�V|�� � /
��p��`�`���ٴ4a����m�/Sj��J�O-$���mxt<�**�]�_�뗜F7�f/$���%pW�kPa��=~�R��6vw&�7ƙ���SY�4S���V�9��<���d�O��YY`�O�ެH[M�a��e83�����_w1�i?����ߙ��Z�T��]
Iapӊ	Ԕ���̄����IX,��'��M�_���ݮ|��$|4�ܴ�/�Q�\=_ưA�%�5��*�?�(�N,?�Q�ŖN���6&�ƲcF�����M�ֳ<�&r�Wm�������v;�&C�L�C���l0��QLǂ7���ЙTnZ9� �-�U�'=�pR�m��OY�l���L�_{8��*�_���a��s~C
g����Zu;d�WcuI�m�fBn�&�����|eK�D$_�u�w�\U6��O+_n_Bݝ����qd���fJ�V�7��s�� vc+`�c`���-t�C��(��y�<b�r܏[� �/[���Ȕ]�c	���tI�����@q�C�N�����N>FQ����OzH���3��"�^Ԗh}�~P�!P�F�H9}�*{t�%���)�ylh�ʨ��&>?��	3��a�_���&�(���tf����1��4{�RR�"�&�LY��/���z�
#��Ke�@���9QC�va�)��~r��٣�2�vf����f�7��㪮?r��m�B�j�*a	Y�_z��Z�yܔ3��М&���̞;6�Ŵ � �"C����|���1l�5L ^C��׻c	ñ�.����/n���(�	�!��b�7ciZ�N�l(O�6}��Y�x��ȥ�/������� ���Ì J�r`��"�v�