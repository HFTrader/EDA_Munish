XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��`A���L��d�>���}���� �3��%���սGū}�}�v�.��m��,���G^J�H_��oɣ �'�S�x��նg�is��}����<��\���*�R�|���co��vg4�5j�(�";�F��Я�o\vE�_�+)1bEW���J�#����F��H]�*����r�����@bX����9J=�%�5�~us�d�Ly��Pu�O�D�!�ɿ���<��ZH$��>��9�=T���#?����a ���aT�(�DvD��J6�2��JꆙEX�K�Κ�0�Ҙ��;J���%l�Y련L�5��+�qY]�r|�Xt�W(A��|�ԗ�N�����A G{��� L�I�f�M!ˍ���@�&�/;z���Ҁ��hCIX�z!R��x
�b۷�rNwe���n�_%Wϻ� f����b@�����ä�2^~���;ƌ�dvN��f���)"�G����5��A��,�w����1��u'3�2{ko�G�#�1�'�JB���������A��+4�uX��΍�w��r"n�x|�H�G��H�E���[~\r/?��ˌ��8��+��@ǋ葫5�vu��c���V[!�����Lr�P`���7A��ͅ˱
��z��L�5�Г^g�6�+�X���@��W���OA�V?0��#�5L����W�Am���tNL<���F�`�3w]6���M���B�ŏ���͓߼R$A�W]!f��<��}8M�BH��Mq����kR��33J�LXlxVHYEB    1e3a     a205�+ڡEUL��lZYõ�������TC�Ei���Cp�������W'�ȫ}�l���X��o_6'��~��-~�T:�n��r�C�k&�R(� ����MN�)7�t-Lu4�`y��\ã�|q�����Ed9S�P¨��K/}�	� AK�~�$h�/\&MDK,����ӛ/җ2�wʜ&�^d��\2��"'��\���eׇi"odPc�gx��"2m���?i�f�k�3Bke�e+����p����'�H��I�q�dZ�1�v�0h˭CB����D"�'�H����d�!�-��<����0,��S���#Sq�R�`몤�B �Ls��[ ��^�1��wbL��Tpo�D�,áx�yJ	Z�2o��"�C�5�P�`f}kci2�=u����2��������~��:���,k�v;J�,��A�z��*�G �	�_��Wc��a�Ђ����.��r�LkE�S��`�?X��iy���Y�"f��Is�����$�����
��p˚�uJ�ר]�BB9Dqd�o��-Da��C����6�S�#)���G��G(w�4&��1�+/��&�7��m|�-D�h�.ч{���k�A<o$ ��N٠B��K_uDt7<x�J�Mf~B����G � h�+x�y���C�}H������<3��݁���K=���`����t�K�B���l��
�������5O�[��b[WЕUu)Cg��x�� [��t��~B!Q���Qt��	
^�ib�ja�t���|m����Η���&�"m�zIJ�w��K�z8UG��ۥ���X��eW{�-��B%���/hƂ��MFK�����Q��[�(�D?��2���ek��$���8�0+�}��"&���+W���qQ���fדc�#!�	�uY�Lܧ�k����_�^ߊ��Vl�uB�`���x����0/ b�Z)�m�`!�A���Umv������@�e���iU��\�3��#��Ȓ���]/G�4Om+�p(�߼eӸ��m��$������ЄY�Ԣ����A��_(�QYo�8�-��>^��y�nԎ�����3ZA�^i�,���Wr�o� ;N�t�2���ߑ*Ct��'9�
��O��U��&`a1W\����b��x��
�d5�h@�bh�~8�����d8l�x	�^��r���Q�^s�k8Vy+��J�]���N�b[S/���1!%�!(���P����)�Æ�A��y$ sѢA9@F��QFلk���qz���V{��_'�X��G͟���{�=�ꕝBR�CzN�F̅�?𐚾%{��j��ڙ|��q�FV�!�})�V�/�7���1�+NQ(I3��|ޗ�y���ӱ����E��J��d��I�'��P��Ɪ��A�\5��a�ߌ��f�e��4����B�K��e�H,��s�T4�����R��IUm����ƛ�>s�o�h[F*�ggF����U [8�>�"����Fg-�Ӷ��6�l���`�BD�}�2�餝+c
κ;舝�6�!��p΍����q�)�.�l�}�&�������t�2�W|%����)���ͦ���4�}������hqN�@!�Ŧ;�E���R�Yo�ℹ"�1�2\;��P�[�����&��<pze��]�|H��K[�+,AVy�`�	o_]���){�R^¬e�=�	Ё_��f��7+�j3)w�$�N֎���؁s�ZUTʦagaHk�ɵ�y�s�=cL�,�dۖ��*�� �z"��G�6�I���?%�p��ՎL��eoa�:��Ø]5Y���� �g`�G����,}�,��P�o������L��ׇ[& Y�҉>~�d֠�f(6�z��G�m#
��5D��|����1(+�ש�������N����[D���b��7�!'=�1�'1iUKHRH2���1!�Z���ʗ�,�)���6�����υx$L̘#�>��\��ӝк��}�կ8Wi�-�	�0d���m��A����:k���z�1���Q�;�P'�W�[F��˭1$����+}�e;2�
�R��A��n` v�{2+U�<,����W�>6�(�p/Y.�����S��W�p��R��g�0t�=W�l�\�� [rܑ����>��em�r��Lb1��8��!#EW��P�\�nހ���.����#���}�y�Y�"���w�%���2����Y�P ^�C�	��@}+�73(�_�����{ ]8ʸ�+�4��o%Nd�8����h)K ���)M�ƛ>�������8S-Â�~w��έa�ۮ�s����w�(F���=���J3gt���T��s`��^�q[`IRT�����#�e�GEZ��406"�}�/�z�+UԂP&�{�j�| Z��n��_��	J�v�Jtzx]S��
x!v7��As�����u�kv��y>�f���2�b,�gEH�-�v-���Օ.�g����
TuF]��g���ι}-q����0!(Fc���i]�i[Q�T�'#��8y�,�8�"�,�E�(>�[�3���r�RFE���0�:#����*