XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{����� �䎃���6���[�[��h�������a��G��f� ��Z��B����`������V�ԊZzw����Z��>r8P̈I=�<��5F��7�"����aK��9ؕ�m�Yo{�w��`x��� ���]n}�N��-\�jᘉ:���z�.�A� ��l� �s�MՙW����8<�o�j�W�|�LTg�/��kT�(�=H��:}q9�qB\��{gq�@;7�4���S˱<���	x�oT�P�3����3��g@Ɇ
���'�mhØY�=��e����IL���08ϣx%$�t�%ҎG���,h@ԏ�Y=0b�obގ�&��&�4�9�9���!p�q0�{P�2{��gD��}:J�9`����ݯ���Vs�˟ a_� ��Hq���ɝ�g����4N���}Ć�r��Q[��cij[�$�B��4�J��ؑ��kn QG�N�W�z�6����?���,'�j��b��Zom���8�J,�j�E��	�����H�@��#6N���*x��[?�]���>�pk(NaE��q�-�wa��CU�o5Ía��8� �}U;K�
oU�je���g��d�n*x�e9�{��� �DSK8	���d�]�;��/���V�]PM��Q�AbӘ���)���"������z�����،����|_
Guxu��@Tt��^*����5�<G�Qek5Fj�&�B9,P�ӷBp�\�-χ�_,�o�XlxVHYEB    2dc6     ae0(�nJ"6���|s����)�+@c����)��'�A	7dMyJ���pѸ�i�Y��'��S�z>t�l�ɏh��9�K^�)�r��&Xb���M��]I,e���6��K�.��u�y��k'���1Ё�
xE|��O8� T �m�+١p����v�b�X�U<�iK�m�}��b��)B�Z�#R�kHt���|�R$�:�XxS��KK�FALc�x3Ϻ��/i�>x���	��jkq�Ҩj��ԣ�M��BuvpT}�W����0�	�dԽTE=p����t����5K���t�g���ͽg��FL�*8}C3��'�30�v�#��dV6��>q�ʤ;�y����jc��P�g5Ț���Q=���יP�ʬ�k�^��� �� ���-���<�R��,ራ)����"1�:�+aH�II�>��/N�v����A��7hy^�.�X�h2�u�V/��sgh$����ol0z����$�z�\�a��b3o��{̈́��c9<��fZ�3�s+|U��R�%�����V=(C��*�����cR���߫סL�0�m՟����7P~����a_�T��R*��4鬲����R��3�W��V�i�����]�oO��Z���%�r<nX@[�S&���G��[��Ȍg£9'�
�4��F�S��+�\�>	��tӘ����*
Yq�����r����Z�c|t$����˛����E��h1p�&� Qߧ����x�R���FЙ�Jņ��)��� �s�k��9[��ۃ��S!A�qJ/����Rq>O�е�DQ���p��B�D/�S�&�6�$�Ζ��n����-���E݋c4f�n
&����ٯ���Ձ�R���� �"A��+�m�
�lp�H�r��vUs��Ұ#(�g�������s�g}�P���jb������:��F�jus�V�9��TM৞ҰY���2k�"!����u���e1S����T��v��Z`��6�4��k��Mg/+��*��;w&�ɇW�}<��|�_�ѕi� �]��ݯg��:+���X?c)eѱ�tH�r�=�YqMd�{��`��j=�k\��& ���_N!9�}�[���Ho����o�\���]�2԰��*g�A84�/��`�N^�`i�)DM.4D��	�p8��BW��e�E��Xh�܍�9ؐ��}�һfl�`���W�uz���I	����	�-����V �xZQ�[���_ajd��l����cPv���ޗ���V��x��]-n�j|D��_l��x�X�d�\TpGI
0?��1������YtW&��| ����%�{�w���������Wp�;Ov�e��vJ�Ig&hm&S?���w[,}�����@�Z�[A�2�e�v�d2�H��s� �6ml_\�l8o��X�����""*Qx�D%m���N���=��>a���Wh�XD i�⩎�1q����4Q�B3�lq��b�)9A��ߜ�i���.�)4��L&Jo�%�Y��0�@��7�������tW ��3?�{��W.��ӓ~�����<J=w_F�L�ク2��[o�d�r�$x�m*Y��ج�k1��fB��	�eC�0X#��Fw˖@�[�/�|�@C� ���[���v-�Cv��x��(�BlO�b����%7�sY�A�c��4Oܼ��09����	_��~��:��=�d2��gZ���c�fg�wo��Aˢ���n�R�-��l������`Pp��(g�%�3l��̰}]���i�v�*�<�jHM}c�͂�s��3^��m��=J�� 'T�æ����Z�7@B����q@��T�j����s�ш�?et�d�[�)[�%�yW\]�>L0��=�3��`�"�-�R�)�U��0ؔE-=t~��V���8P�L�[�v�!�yV(�qeŘ!�x �~?#���^)��K9�NE�Ss��Yl�c��ʃ��a���yt-5��4�ls�˶Y�qBS� ��Q��y��X(�n^��c���A\�:���'�J@0��h�С�H�6S;���5�M/�QM>��y�ڽrTf�?[2�@�y�'y�K'�,�o�ĥ���㘏r(U�gZx05��6�޻�q�"ּ�"U���n�w�l�^��;
{�8��`?*k�[N�}3�]Y�v�?�9H7��b`[�`�������5G1yҦ��w<���#��cEbp�tU��ys¦���,#����������1�[��]���xu<p�)i�ϖt��@��]@�VN6k�we��݃�����x<� 4�̜<�ˍ''���ߌz��b�|`�6�Hp�QIҁ��$������N��@Ѵ����Cp��<�%5U�2���mK���#T���ǂ�%��(7[$7���X�D�<��(�3H�-Ivu�\6#��$�ky��<Iq��#a��\������U���pQµ��S����Z�0���z�<pۢHx�dN\A�@����%�Bp�X�7�x>H�3����v������tI�] ��xJ��tā� ������
b�'�^{�A�d����"�Xԇ�b�[�\��C�4��а���o��ڈ�f}��t��#N/�T<iy!&`S�����}���ߠn�&��um��@V�=�@��Pl�9�i�Gp�b��K�#�CE�r:x0E���aTt��ǵݤ$������5����@��y)2#8.ce7a�����L���,E�V�N