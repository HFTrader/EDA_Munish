XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������
�g-Pc�qY?2}�զ��	>�M�Ҧ�`�fBe��\׀����;Cu�S�W�1�� & ݞ�O��O��\���m�-v0�<��
��ˮ+�t��Ro��Y-��X T�	�X�d�~�|
fe�Ъ�v�	ġ.�g��|���`���FQ���~�X�)�	��MM��[��9�KC�Ʃ&xw�5�+��Dy˱�|�6��/S^�� �P46_˖��݆$V����ض�Qεz�����? ��5|�Z����ˡ���Ɠ�A�4���y�f-E����B�i �/�yw��k�,��_�K|�w�9t1!Y}�`sY"�|�2��3�1���1�#���}z����K�� ��Ո핀���>M���������8Zw��]��TD}��*+V����;��byz������R1���+
� �7����9�|�����:�t�(qF]��J6�<w�Їr5���A���b�A��{�I	�py��kXw`>��V����t_��?�t����a�<����҇�!N����*
"���ݫ5 ��n1o�I3c�6���R�m�8'v�CC�#Ry�R݅�E�XR�|���[~��ц����_GWg�G񬭴3�h<�x�'�lA����3��S����u�KK����zxT��������Ҡ���>,g���S�\��D"1���G�Σ"�Ӛh����V�p�~Y H�'�����︣���Z\��#��XlxVHYEB    9efe    1be0p�*m�G{�%c�R�٣#�j�1)4	^̀o3z�u���C����6�ujL�0n����J޽ �x_��i�y��~���p���|�8�z���y$f5h��c���H>�s^-�RbZ2�AV_�	F3l��'۸Wj�At�6A�X�M_�b�Zl�����[|~+b<��}�����aT��.�j<m��V��ԮJ{$&�O��W������\�ʸY,�����*�x�g1����jբRt�³�b|]<�����
n�R���� J�z��yU��m9
;M��+���t�,%s#\��?!���	ܤ�^p"U@�bB6���*#�x_r"@�*%���l�[]��!-󐤦6��Dŀ�3�aQ>L��[Z�{$w�����:[;1�
�[k�������κdƇ������-d���M.cL�LV &̣�r�kٮ�m(v"1 ���FA��82��׺퉱a��i�Z�&I��X�tv�/wP���djR�IB�����h��~E��l�v���0#'��^����6�9h����M��һ�5�X����F3��|S����f�D��3R�n�'@ӻk��.����&��E�cZB�ց��.�g��5�������5n�I�g�i�vO�܍Eg��(0��Yc�?�g��͚�>f��QLR�g{ٕ)pq�up��")��䕂�H}�[Y3BAaZ�y?`�EǭH-<�X���_&�<�&:����B��(,�aЈ��:Z�$�5���A[F.~�w�c˖;$b��`�|��6[B�M�?jes��S�0zD�Bq�~�M�T�Q.:|�QzE$P����\e;:�5�V���T4U�,������S'U�⍐i`����F�U�wbgk#m"����'�_��n��9�����
�ƺ�l��ߞ�$>u�8ߨ*�:C��ѡ�;��J������^�C��� [��4%�ʩ��ч�H���u�_�a��N���;�!83¾|3��\�WH�z�X*(A��q�z�C��i��I+b����g_.�^�����,�@ ��2�=�B��Q�0΀d����=A�ã�4��5�C�X\[��ՋqG�D|�(�w�қE��7�]��������4V�L����w�Z�#n�*�ZS@PA�	8�P��X�Ĵ7fF��s"��J�+A��)�������L�*}�; mƐ��jk�O]x��d�q�a��4nM���)���rh����c!]�Ή~��z�i�����������邹Rj�hs��N�٢x�r��m�-F|��π�zW�EY��A-n���KW�:6��0�!��L���+�����^�������t/E2�ת�-A��C��`�S����@��b�Y��čωk���φ����f�|����p��L5�#�ɵp��6����1��ݚ��k�f����*|�ZR��㺥sr'N+2$����KO�	 �n?r�ԇ�^�������p�!J�dF[�fq(ȢP���=Fe�L����!*F���\R��em��'~v�v��%�Z�0�0�ݛ�$���"��x��?�Wc�b�5��CR+Q���7�����ݝ�<�� �ػ����b=�q@8�P�Q-�t*ϕ���LÆ4�AzK��� s���|��3r]��+ce�t^t9rHOF�����@;�|��}�b�����>5D.R�Ư�����7�ж�p�Q	�PbD@Xx><r���W0)����_i������¢��&���ā\����� �@vF����;XLP8��	b�!��Lb/�Y
�yW���~��y���B���Q���!_�fJ3L��K�Ŧ����~�h�S�F�_~!~�A��D�K�Q�(Qr]�F�2��fYP���s����*O�NJTP��T0^� l��j���^wa-�+.߱5�0�����%4xѿS����3�yX������-r��̏Ы�Y,�غ�y�N��ȈWȆn�9�XF�����"��c;,![A�?�c\h71|>��p�y�б��	��|j�{	}�'i[���{C�@`�a�.�Op~��$���ʏ+�Fc��J��ˈ���y���ݍA��I�Y^�~Y6��Xa��: �@R��r�?;���/�2��Q&���tbw��d�����nsz��{��=�cH����F)��$D�{&��L+l���q��x�2.�Fҝl�(���~w��w�.��-��9F<b�D��
���{��>4M���8�8�R��B��s l����bS�X~ݫ�H����9�\�о�U�C�f�(�FuR
gH׭�L6*�R�"�(���yWy��9_�r#�������*�.e��	>F���]$n���ݛ?�p�Y���=�'e��{�/m�k��^�1B|>�1 #QSl�R�䷥	ki��Ѻ�?'E��m`%#�TsW�X:������O>��U�n��0AT^G��B�(�i�#��m��c�^������I�J:/�=L��iv�D��zR��i|pD��(fsWU�M��'�L0Hߟ��H��/ƕ_$0�v�������C3��ZϺ��G��{�dw:pUg�+���u_�ua-�9m���yxŝFݔ�	��� ��'�gTM6g�tV��*z I�,@͈�O+�P@��_���%H��T�8��}d��.q����ȃ7Tb�v'��GΉ��'�)�1�Dl�81�G;�͙۫��՝Iwʟ _`J1y�+N���M\��M-��X�-�d�	��}��Cd��
������Z0�����^�o�t@p��s�ȹHN�Nv�2��:�m¦�[��6���^�^�6�\/�Ö��ެd�����W�A�4��j�������ff�FF�Rm5�w�I����A�d;�uR_F��4<�(sPB�H̋���$��7�h|��Ş~EN�����9��/�?<}H���)���) �O�{W�rµ?�n����p�ǊFrZ;C����{������G�쯩�W]<o7b�xb�Y�+u�����g��?�+�G���+�.��c�t�ԋ@��l��`�0��j�Q�h����N�|�?��ߋB~���x��C��mp�����爫�|�LH�M�B5�~��b��y���g+y����FL��^op�q�.-~~9B��I�n1���G�C����U����ٷ�T�}8��˝�9j��GyNV�@��C:��_%7�	 �3���`�T����	�S�1�LDdŉ����|�v
H�I�m� n<郚q^^BF���0@I=�V��}�����Ύj��~���T]T���C�y�J�1��s���hSs���-�I�&.�=#3�����@�{_�xO:�C������������ �\(���n	}X;;o)c2(�-j��o	�92O��ٌ�� \��O(�ȴ�C�T� ��ܵ���r���o9!	Be� �:7x��<&��ʑ�.��S��������ݓ�(��ˢo�Q�I}W�xngk,�+��3R�Ƈ7��R8�U�XH�Θ>���ln�*�^���|q��#;J�5�3����HO�'���@����	g9�C��}��6�V|��S"��	O�{��*޺l��<��?��9���RBO�6��E�A7�QІ���Vׇҧ�q	��dfg ��R W�)����׵�[a�������l��L�)X6���֪K��|t��0�9оN�YA��=S�?.���t%է�|�yS�Y|�蝒��4j�9���#��ϑ0m=ש�/[*���4w0�N�6������Z�U}AC�������{m�Ķ�~�\{�mGE'
�f����<w'� ��Y��V#�z���b�����j�4u7�G>6���]�c�K<CR���% E B�m�`���g���v�k��"���ji�%�ɳbR���?��*ؽn�:�2��a]�I��5��t�� ��������������R���=u Η	��R��3���aՒ�ʽ��	O^��#�xD:������Z�E�����Z��T������$^Rm��'\RQ��A���#(��MB�1�	�%��)���@���{hk0����1��o���qҲ�G�{��VB���=FX8E	��{�	�=3J�jz�0�RS �p��[��@'���;�j��۩���1�A�}{�1�U��Pz]����'v�c�q���2�2ū��T�a����!\�/+�AˤsQv�n���0�n�7%;���g��;"r���J��K�(r���]6p��Y��C�K-�6J��$ܛU��I;�M�?UCso�!a;��=%xkč%�] ��S�eȯ�����v]���C�3h� [����헋����2>/���L��������(�x!IQ���f��*�X���	���,>�l��=J4��
��νl�E],Jμ�2�Wb�q/��IH�R��gb�_��|��4�05
8NF[�,,�S�A谀Wn�uzĶ"j+�rn���>i�{�%�b/�eu  9���Ԭ�c�d��\�I5׬�0��7_��)
%kt�d�uM�>�I���.���,BAf�fAx=:�`Q�_6,Z�&�馱��R9<{�p)6(L��Q���^ֹ���V�>7P�؆��aC������B	:a�e�n�Q9|Q�ų�d'^��mr2EiE,�쭇��ߏE�MK������P%�c	��'�b�
-���n>R�
ѱ۟��Y�x���r�xwT�Bb<�y�2��l�tĻΩ��:Sᗷ��H)��#�[�zf�pч��|9<Y�
}兦+ܰ@/�H��*������t���X�hoK�-�1NO�`��:��g.K'���������n�Z�2D�ĘEnJRzqw���)B�݇ۦ��N�DV��`:1��ȏp�:<c���o�kN��Ss�v�)������5��zw2<$��I�b��7�ʍ���&�lp�汆_�Y�3���V8#����X�]t�"P!x�.$���(]��筠�%���&�.uI�_�O{�'\U^.��x]�\���C�E���̣�w�<�Y>"ű�ԕ�� �a��Q�paEn!����5ji=�,dh�\ʻ�O�ԭl��
�Ƴg[�~�!c���_�6-΄W��+,ןhq�>~�V��[M o�B$χ"-Է���i/�0�Tk�Ę�)G�c$E��$�COy}Z�m�T��\-�e��o-�C�o��2^�q���e���&�`<oWgS����9��PB��1�a��/��n���ۓ���v��M�^�n(5���dAZ3N+��i%����Ү��w��������u���������!�^gEQ���O.��RM�_���~� D>�T��-�qvܓ���2��#�t��AR���J ���%�T[���~�q����%�-:��0��"i��cQ�� �����	h?�R)[[�ah���w<\!��m����pH�g�n����I�+�� �h�� ]Q�������2Dr1\� ��bG�!J������Xl]��Ad2÷^����d\3|��������G�N�c�䆹�C�0G�g��WyJ���fH�p?�3(� �$���@r�WX��;(�cH9�q���a��0�'��7�
`C�Y�?-��5��T�f�
T�	�J��QqZ�p9Z�������w����5��oA�0�?��g�%��PN��Xf��׫9!�X?�xm�s���hv�����Ђ�B3�g[��B�î]��&���C]dr�Zo�}�'������Y�$;؁Lێjf
�Q?J�s7ɭc��@�ߛ�&�-Q�b���k�f�$܄���`�rEByoQ��B�=��f6DJ[�^P2k����]L��Q8�>Jv�v�N����� �Z��bu�I��"e�⼵�0���>�y��{%��s�,���{��?���]ӳż bY�+o&���螗g?�K�n�p��+���	i\��:��}}HR>�t��SV�(Ϻ���t/�դJ\`���B��F�h�} R�����;�F�/�V���4�u�pM��YY�_د/j��h��Ǫ�=?N�����ՌA >�%�g�J�g�#��=�o���(��k��<��|�pƷ>��)�w��ξ�f+���<�BI�aX\�ZT�K3��E_G���)Yp2�@a�S!����l�&9�лE!+�N$�v\��Yg"δU�߆s8Aq�3�be������ZF?�"���G,�ڬj(q� l�l��[�#���<��6o(��'I�3��XD�GBLU�&��e��nLlHߖ�W1��=����߫��D��:�NKk�������7��}�*����������+�Q+�r�k��'�
�<.e��S��u�\|���?�$7�\�y��_(ױG�֫.h)e�G�Ss(��&�uA�7voл�ب�a�+�P��a��Hf��Ê�\���硍WY�g��r7�y�.�rk�����@��t��7�C��f[Y`qC@>g=��D�MF�`�L��qL8�8 B��=A�ߌz1��z�?fU|?�SB�8#������q���
��8�\�B�~Ǝ�b���á�՟�����y[̞�FC�15�&q�G��b3��{��ߋ��z���b�t|t2J@-����Y��K4�^�U,U�)5�2@�ְ�?��.P�&�Jx�J�0�ܾ�VG�uR�	���-�>
��������HLݱ��01���|�*�H,�V������'`��&���5���H��	��+�`�oh���Y%��7 yd���D�c=��+�fc�A]X��	+ɞ�%��NS��A�j׻<�n5��Ⱥ��7�\z����}.HAD�d���>��]�k^y"C�],�Xv��q���Ƅ�}��q��P1%���{���Ȥ��j-^sK��ĉQ�߄���c�@F���λ\	D�5h�y:�$�6E�@���n�w�Ua����?~E���O��̮]��Sp�S�0~8�ӡ̳�X��R