XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5�IT��3������P�[�Q��d����2�f/�l��j�M�x�\M�!2�AF4ط<1����p�h*����`L�ht�	�3���m�k��+�`|)�hZ���0��SE4�
�Օ��2��+��*Z���5q%D������FweI��
�ȩ�	Lm��} ����79g�'�,
�Z
1N���o�Pqה�[�4[v6v�O���,W_��^��GQx��!v��w�f�k���h�Z�ğK�K`��cP��;\�^�R]&�hd׀
����ǲ^#�_��t�JC��D=߯WS幇{�KS�0�M���Eq	OQ�֗=km/a�r�:�oD���i�s��U���g���n���*�夂8-�E!������WFҤH�Id����k���*��9�� pk�|
q鑩�|����A��f�V
��a]:��YT<��0��C��-l���_��e.:it���-�,������g>�
\-y磫�~��H#�_����
�G�[&�m ��/�C\��S�A��=#M\��q9$��s�#��Q�rM*�QX����4�wp�T9�PpѢA�Ͻg�(͓��/��N�i�e�)�y����0��	�UH��z�����Z-��T�����8���@�`��-��\�u��=�>u�hs�h��
m��=fd���!a"~'�a���A|��栟X6%������<t�RW�r�������挸A��4��ܕ�@+o]�&u8���7�3�ku�o��u8��<!�[XlxVHYEB    1959     920�#�;A�����0X����<8%�ے)���Fw���v�B�ܘ�xOr�j�X����Ώq_��~A#˷��ӱysC�L�G4=�hr&o����C7
4]�-_�^��LS���#Y�iIX�fFh�����.BW�����q�Žj�P�H1�����91��I�_݄���͑���5�uNiy0����q7R��pH �\[�07A �}c�e�)��� Ԡ��+�N	�Ҿ����}�}�8E�e[���[<"&��\���T{���y�����=�<���z�kR�k&D�2�S�God�m��O�2]���Z�-��"�:��KOw7?a�iҏ�ڤ�I�@]�y�	� z����rP��ש�9���w�X�=��'rl�[0�.�4�q>P9멈hǐ����F"�(5���Ѭ�~Ω�LUR�+U���Rٔ�7�t����CO��2���B�
�N�m��5�{`\*�Ӵ"� �M�y2M�O3�E�_J�i|x�RG�$W��9��+x��`f��ۍ3Tj��:�g*�XW9����7	Ê��Rѳ�+��Ȥ���~eY�1@� i��8�Ñ��?��{����mR�vt���Zc��;��V̂:�?<%ʈ��n�?��G�f�]Y(��A�a�>���U�T��	��� �nd��{eV����}���D.����۲v�����HIb׺����=�����@�`�))�>���E�&`���s�+U��RD)�T���:O�`�E7��h�t��t
~��E�o�7 Q�TT�P#�4!gz
�r�٩�0�e�\�;�?�&:��c�x������o#E�۳.���m��ʨ`x]��se�O�Y �rȆ%�u��Z��A�L�0�o���~��x�dʴ�S�70��v6�5��J�D,�ǎc�9im�G7���2a�K-H^���݊��C��CW!���-���k��8NAH���*��֦�M����$��e�1�*v�a�cv�P=Y���u��9U	��z¾0+�f>��<���H�d�B�� ,p�f#ǚZѻ`\ז��%��R�DYV�?�%��><c�eh�]����/�O�?gim7u��EЊzI��252%�Tz�?+�����s�\f�����*xB��H�=�S,ٿ�*]�6`�i��]*��a�}<=��m�W��3�zz��fl�rQMRG~zɻE?����>���z6r��n$������`�3��>ȕ���c\��u�:�ᱴ���>po�r.�/��i��,#j�(�`tv`E(N$�"A?�v��|���wa2��gqx���/�#޺����_	
jv�Z|���� Oz��|��B!���ɭLp=������b�K��Ag�*�2{���ù�&�������l��X�%��xB���h�ڰ<>����H��0�V�i@������G7c'L�K8'Z�|̰u}��5u�)���p��ܝ��o ������0w$e%ޏ���Q���el>�-���(��OU�A$b�`�m�b�(�`����FG �O�l�d)@o��S[��������S{�w��@ϠK��~:F���_l�_ /����g�s-7��r���0�q��%KT2��X
XK<4���/�CD.n���9-�dv���S�=p�7��%|�jj���nn{>n��w4p|�,L�����U_o�c$K�
Q]�?�M�ŽUiO��?�P[	/���df��J{a���m�^��I���jj���X��1���*!b��v��IF�i�����H;��9`�L�#���Y����mS4���[Gf��ix���n$}�or���X�V*4s�
���3��*m�M��q·�_����m ��Z�W�\�s�OJr�P^�@3�yef���v}V\�Й��ǰ�oJ<m�6ҹ��<Fo�A{�F��;2�FK���x�v�_���# �Y&ֵ[��β�ox�S-�\�3�c�rv��������>��ϕ�:�W�8@2ov�ڡ�-�!��GD	�σb�jZ�O�r���Gѡ�o�?�B)�K��2�=�. �(�ˈtf�ھ�O��jK���O��NGh����^)�,}Y�ӿ���Zyqj�CDD|FjZ��K /�Ng���]�ҵM+i�'�Wm����<F���4	=�4_����Ѹ�7�C�$�A09W�1of�!�@�X(��VnXѾ6���x�g�G���=-o����؉Ǡz�8�
u�����H�����~��������?��������|�o$�d6Q����i���dR暅�$}��,�$�S��v;����y�&]צ�c7��$�ʆ\$�g�6������٩	�u�i