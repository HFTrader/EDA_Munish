XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����!�k^��33�B�I��>�F\�.�%)����U�H��L�+g���UWf`A���>��pV�<BPvf�[�2��)��mѫ���]	�[�4`�,Aa���b�CJЋ���E�<ބ�o����.'Ð�R�#��55��8�5��,��=�d$�n"��pi\PC�Gg���4��9R{�7Q�k�[���T�b�a�nZ1��Q`����W[�+^��޼ɱC���7����j��I���<��5Q�I@��K��������q�S�!��	�OM��9�5��
�����*��>���]�?�N���`��j8��Z��aL-��\�\9�I�����^d�X�]<R*0��0���mU��e�?q6�EJ�,��Byf�c��ЗRwmL�J<i�k���@�v}݋�՞*�o&X�t9���ڦ���B��sS$c����Ӻ���6��;e��z��l"��Bv`'�ADJ��|�n3����]��U$��ln�&�3E�}��(딨n��+�2o���f�{1:��5��G����׏J���*���Z�_�m�77xU����QҭS���A[1�[I3��UL>�&g]Yr��f	�E��a��A��V_t�x�YG�ÌN|h:�h@�u������a@/�;Y���i��b3���>̀㓬��{�{̘x��x�٫�+;KC�W[p��$��J��c��trK�M%(����;5���f�X����$UKy<!�uЈ0�V���pA�:QV���#
��[@d�ױ��ݍBXlxVHYEB    248e     9f0�p_5y��jZ	�:����47�x��6����6S��G��~��*w^ܥ#�G�s�B�+rs��f��}�2p���\�=!����8Wę��?�[j��,GcT�6VPd����ѵAP�d2w�ʓ��1�Ε1�?���O�`p���9aԓ.a�ф���xDz%�u5o*�ѣu�M���v8 �`)V�ZNd���J�&7��F�W�G�����2���������V�y_x��f.@���"e�Q% ��\C}��l����]Dߘ�s��%XoŸތħ�|���l[�q��U�e�?�k�ʉ(ӹm�֮
pY_��F��ܺ�1��ĢX�ܧI��K��ň]X�����KK-�����W���YW�!����J�3t*K�
	5_w�PA��.r����1O`��\hq/%����u-V��'�ñ2�lm���ws�C�>�*r&���İ�N�-�&Ii�K¸���Ѡ\��ɿ1f��;M���-c1��Eã52��|�g�<E0d�����@%��	��v�_��d�nc�D��?.�~�z�4��K�M�\Զ��R	'Ⱥŕ�����dk	�꯷�#��[�L	6XuVP,��	������~r旮�p�0�K�~�uT�fӹ1��t�
h���\	���|�����i卒l���IU$ݍ���_�0)X�O$���� BѬ��(�&��_l�I�������s	36n^��4����n�d5�ܛ�Q�q�b3�I��܀.��AO�Q�J|�eH/[r����Ҭ��jA��נ�"i��4�0�8n��$�ߩ�0Ŭv��2"��̯�)�J�^�O���X'�l�&l�.�B�J��b�-wE�e�6��ȕK[��gm�O'`�v-��ƶ�̏��+%�φ�A>�s<�r_��#X>�%q��}3���L4�3<�ZG�?��t#�����\�O�tr��T�{���t�2��U*/����%�k2� `�m���{���.к����������K�\��=�ڱ��H�l���Hl�*���AW���$��M�ǽ"��:{���������=���"������l{�wez���+�ZJ\tNR��JR��{ɴ������Y"����V�Xb��,
��GQ�[P�H�mA�3��(��:��f(��~U[KA����bu����a?ř����i��>�+h�7ǳ�{�^�����#�ώ�#�7�Z�~ �g}1Q/$�Zc\a-IPS��� 	�-{��Yj�������ޘ<M�%?Ւ� zgܪ5ܓ1�^*��@��E�X��Q,� �,�<7�]���~]3�����^��5J�~�z�y
�L���b�	��i��Kq;tl����8G�S�-��H;�T�60	t���C������\d�P�Pm�^�C� Xs'<��g�� ��F�b�h���[�J��Y4l�R�1%��3��\	�M@P�%��Ě>5[k���y���[��]�����������PKtQ���!u<$�"	�>�\��W�� {V��NΥ�Y�d��$@�`ķ��`^&l�Qa�.8�<�"��ᕨH���$�ӑ�G-6������T]\�iށ6�Ǵ,]�����[�q����$��(��'<;�q�嚘�TKr���YxUG~�oAkB��
�e� �ș�n�W���,��|q��L�?9(O��iYN���:���:)�]��	t�Oʮ���$�^ ��̚ljI���zz�_��gf=����=Va�l܇'3A`��Z�d%𤱣���չ�u�hg�zM}���+��}��d�����߄a)�#&�j|X-#H8�'9�<�iC�C�0���u��ǔ���&P�9fN��� �G��KE�Wz'�c\f�ʩ���8h
]6�y�T�� ����;d�I%t��@��xT���'����U���a��9�&�f�@`�c�.�|�v�U�z�0;2���Y-�O=�H�+ �<�
03,�5�j!$븇�[��D�g�oU5���{�6���/���*��e5|o���d'1�URQ��z��eJ��	����쏖X됶�s�At9(�>�^�R(�>���: *J�v(�L�O(X?�#$z��L��Q��)�O�����6';Y�!M��ʲ�gO�x�M��an�ڮ��!z���>��Fv�G�7�	�d���#ǛAm�q���n������f~T�� ��d\П$�
z��u-Ph�>�8�X�@�L^�@wa�TI+��i�P�\ Qؒ�������=zi�+@i�3��o<�)
)$_����yo8J��-���Ô4��<�06P.m�0*�wܑ$��,�=�4��Ȧh	�4��-�)����91�A�:7��"�4+A"���I�A�)&��%tb5�&��1��YEi+㟚� ۏ��A7����+�ױM{�|���%�k - #.3=��Z��P��0�>vy�k%��vמ�ps7��O�&7���lѴu�
ܣ������
W\o�4���+6H�)7��J�$�