XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����>���6���Iy�#,�[	��N�A㼨�N��}�ȝ'C����-,0\��t}���������ζ(�oȢ乶����2`��r#$w�j�F��wP�t+��^,hN0�p+�,�"�#D0O���i�R#��B]��Ҍ�o�[U.q����)��˔�[�' �X��R��I���ݜ�[�e�Fgo4�,��)�ޔ/�s ׁ�eT�ē;���1�/ґ1昪w��en��D�⠄S�Q�]λ��]8�PQ������ć%�yK��ӌy���s'0-D���ƙ�%��1*�V=ĩv.���`�V���xw��Z�Eg��i�U�K�y��p��~�+��Ho��,Q�uG�M��5�=�ƞ��I[gڦ���'N�/�;B�Φ����&H���;���тZ{��`�9��7΄U�;��{a8=��}��r�Ώ���:[wٍ��g�J� r���|l| ��d��W�<��[L'� �`�
;5� bq�doP@I6���S��: И�f���_(a���F����S��p�{�D�](�`�+⺬��$�c)���̹ڝ|�=o���E�Z�ޮ��2v�Wg�Z��~��Q"Έ�G�J��/X�l����=�$]IP���ɯ�lP���3M�J�E�m�-a�ܷN���������j:\�3��q���j'=��uce[Iݭ�j��G�'���`q������	?�[m�����0Yx(�ϔhXz�}v``y��M�XlxVHYEB    4f43     f90�Ydq�� ��2�ğC�@+��E�BPM��c���Fu�3?����>��o%�u��d�xͱ�4:x��lj~a��78"�j��º7Q./����s��[ۜ(R"��6��*��(%����8�F]���~�MS��e��fR
���Jk52���#�~Y!0�@���ȳ�����ݛ��ro|j�0�+ SƬj�`?���P�"��'��	X�O/
����USt��&��J�fBk�DI-����U[�� O���1�b�5���|�v�Ѷo�?��/c��݅|�{"�~����3�O�\�t��2�Z���7[β��m�gu��g�u�q��2��0����ۂ�!n.hQ
�_����gF)���T��P�V�GcH�:u��f>I�Wh-�/���}.O�V��D_�8�
����<>$��#����w��A�A�\Ⱦ�.O���q��1p<�Ȭ����"��4�ԶN�}1h�5t`?����w�U�>���a�%�'�4)�P����A��W�;I��ㅪQqڐ;�&���������ށ�����H��݊[�H:`n�b�Z!�z���Ae5h���aW�Gq�N�JMm.��_�g�jk�*�.���J"I���G��p�y�{�vU���?�<�C���u���R?'#��b���WPc��pp����{����m�L�\^V|Z�kE�ǉN�R�bݳ0���VOK�
��r/�e��,�F�����+��e�yu�7lK:-;�
P��~���/�y�s��"߼�r���]�!����;�k-ଯC(1�FӋ#��	��\�[�������K�Bz?}�\mD;��r�{�*#OO�V�>����q.���*�@� ��4�.��|�o��������a�I���b��G�xȠDZ��_X�u?b��	!�4�G���ûq��Ƒ� ;����<���7}Z�(�_X��ܪ��o�kNϑÖL�̾����͠>v׉$��Y����c����eZ����'�ۖ��Ln3:PB�͍,�k�5t}];v	pR]�#4�YGTTm����t{tR4�ױ{<4���:��Z�O�Vi��{�N����qD�����e�k���P� Bn[wa<
��6�RґĖ��c~3��֙XyA�ϛ:~�="*�vG�:p�h�&�U��o����r�|��f�z��:CJ'�O�[~q<���!B�����j��3�0b(�����#�k%����_�)��B<�ښQ���+O��S�$�/O�@wG�T2drSO�V�w\�|����������p��?�@�Q�\��Kn���ǥ:�g�>)W(��q�3a�~a��Q��T���İ��_Iޟ+l���ᒇˁ�ZR'�W-�����/턃�<ǉ�1Bλ�+�,:8L��M`�^�������A�$%q���R������	%^�A&v��%.�52Ns����3F�T3������'�l����L�������²FÃC���,�lq� ��x��#D-��V���L�^*�p���M�ߩyU[��w�+����,�rJ,����Ƅ�yA�r�m�����=\% cl.�c�^/N��]�CHܻV�1��F�80+�=ߜ�q�C�4������8��/v�U�4�IΛ�s!醓���cvg����Xtifq��xjH�S̃Q~���bG���\n{���-�i.�?{�yQo�67�N�*��x�從��,U�a��}d���*�-Qfߘ��A��������5�k�5埪�2��olRIdM�B�ΐ<.�Qj�Ԙ{r5K�������'N;�\��{�xхL^;Zp^:8�ż�AS.8���(d>ɠ#k~�.o��5����4�6Qt9�yK�c����n
����8�U���ך"dP3'�s��uU���u~��v�	�V�Z��U��8�s�m�O����/�Y��6[�&�^����U�4bCM"��6.�3�
�sC����B���pۣK�}6O��S��V���:^NA�~��ċ�W��Wwәg%?>��e�cjQ�k?S�2cX���=+��:���Ňz��ғL@7��>0,����i�k��p=q�?�m���M��lw���f����L:�t��L����-UXrx�rl�Ϭ������uӰo�<�7����8Q�CSp=��Z�hz��}�%���[��Y�j�R��]R0ҥ�fH�է�-�?���@j���S�wG��=�G9��y�.>��A�1��;:9-	��~"]���M�:���P�BPؗ�;��ԝ���7��Eͭ�,8h��~��n���(��Z����+a���S�C�]�G e^�\{im��V����k�e	�[B��A0�1T{�#{������T�;������]�	��k4�%
�����u
������1�lRtA�PA�~�t�6D���DhY�I�U�Y�`t�u����6���A��1����n��Ў�(6BD��<��R�j�4`�A�ߛw�f�L���m��a0�z�r:4e����<�u[����x[z�FU�V]
�Tf����v�:ب03Q�@�d�:@U�4{֬1�Q�#LF�C�>�Cr�4bw{��Ԡ�!R�+]���
��1����!�w��n䣹g.�%2��e�6���?���Ze�V�3��T�uQ�������0�ȟ�p��� L$n����+�b�Y�Uƚ�8���B,���w��k+[���Rd�2�
{�O.����xK	�S@�"?f������',���j����1p�ϭo��Xif�R��371��k[�/�[�f?�+��m�O��A���i��
�DO���E�BG��c?������63�AR��^c�'��$����@�As�l�������8�>nN.��@�W�Q��j���b.�ڵf0ݵ�01d���H/�R�CS�-��~�,�<ĘT�je��s$	��i��d�O>$�r!�!�EZ]�끣p�  ����oީ��,��^Ӂ<2q:%+JCX ��8�+(�E���W�%�Qr֦��L+���05^��?ɆEd�D����`�a&�F=q@�b��^����n��FǙ����d߬B13�r2���drWE�͚���G�N�ߠ��&$߽����{'�(֙�"7&:0�0������-a
"'W��6�2��J!GO���b�ũ�ԍ/�1SX�j��7C7��쫴�k������&��6�o�]$�_��}G*��v�z<�r6�{z�x��2���Z���W�%�4��`��^IH�w��bc����Q���P2��'�xp1�A���c�6�mZ��'0m��"Y>�H��Ɠ&�
xPO ��
�ū�u3��aE�`�r��=�En�&,;���=z��f�$��d:q�+�t`����*��S���"KQ�!>�R5�耵
3����.�����Gӭ�g:���6~�yA��F�l?�	���$�#R�4P�b�7H�/}��L��'�I`%y23+��EY(Aƅ������eܷ��5�d-��1���6�T�
�zH�E�K��u��A�!�_&�VJ
XC@nc����C�A{�h,�3kx��D dF5�E�~��Kl���ntMYF�;�e~9�4��Me��N=�j��O�;�c��T�� �ezܭ�wt:��'4�O��1��/�3JC�=d�\��a��;&�3{�1�?o��J�՜R�xo���Q�7ENY����"�Hldm4���#)�B��K�|8)�&���'����EA�R�}�|p�)��H������C��(�tz|{�u��I��uЗ"aғ²��3rO��l5��+��Ο��S�����k�yn+T岂T�:��T�Y11�S�K��9��+