XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��xx�}�k�l�T��*\��y��	C�.#Z���:�|U���nI(y������;v��� �qS_q� ���, ��Ml;Ce&���Cp&��O<�5q9���s�B�³�M4����Z!Ę,�%;
�h�.�wk��w\���ލkBd�^;���z����>��Qc"Z��n��!i�x�p��� �+�=?�����&�#���6�_����0�%�4�'L?�k�T:'�QБ����~��d�9}/~�3F`�#� (^?|�R�����%�_�ɟ{��J��I�E��<B�jN���� ^]`��,���`8�K���W'_[�*��h�8��$���VSP5�e��k����f���S��I)�& ,��.C� (��2+Q����X��1�rA�o�MKc^p�ϩ(Þ"���з�J�9�:-`��T�ß�ʁt�]��x����B�g-�0LM%(���nX�c"�.�
�/#>�Ѱ�|BɅ��w82H�V���޽z6�q�����9_�P+P���4�����F���ʩi�rk���X�`��vµ)���K&�z(�2���O��ٱL�WMmJ���J�]�P;7d�`���ۺ�J��Bmֈ'OL���M�y�����H���A���!0$X���䨊Q��'I
,[,"�}���r�o��f�
�>�dI-Nov7b�{=��t�o~>Ɋq[F��v��A�$(XlxVHYEB    9de1    1670F�d���I�C�1�*����G
��8�:Єn���V*) �\ց5���u "��^�o�	�ǘ0�a���ٜ�`=�O<�p4ű�T_��raWɵ/-��E��XC:�u��Bi�I%X�KTelh ��'ڔ�
�����9��I�湭AO#I���f��7�������P�������I���%�<���M���ǃ���6�go��pߧ��
�ڍ4�L$�ҷ@�D(t��կ�2�r[�u�(��y'XBF�	wm*���BG+)���_����76w��d���&����up�x�)�h��{U�d�x��p�u��N�M�  c�RN����&���]���C��m?�Ǧ�c#N|
��O��V�9�� &Da�ax���
�}%`֐d䵳D�6��ZM��i�50ӊ��"D%��Nx!%�d�S���rDI�Ƌ�����2J7*�(~���2�����V�ཝ!H��k}���ɉ�t+��q��+a��1�8]�+<8�z���hr2'7@*3z"�N�b�XD�9
���D'�M�z����n*FTۑ���#S��T�q�W'ق�_+���Ջ�P�9���fk�fH�������8����?�έ!��W�o�(4��z5��A����+�*}&.\�v�ˎi6,�'��n'82�4�S�5v��˨��=���*�f�Ua]u�y7�9�`�8���֕z���B��/�z���;X��~�]LȀv��_�����(]����(m�	��v}���7r�Vf�8��j�ԟ�)���g�̖"⏸b�����̴�f�-chz`+랇ח�ߊ}vY���fx�l�G�.��,�r$�#
�@��ꄨM
c-,d��U�$��kݟ4(�O'�8�Ƿm<ج���m"o��r�\#�7�MU��t��ܐ������@d��xg�პ]���kc�t_`:�����`lp#0��?�UT��KPE0�a|��퇋�-���>�iЩ�0�jy9�r��x1�iU����
a0�B�cf!���;i_'A3P������4��m��J8��^=���a��G����\M���pߎ��D�Ԏ��m5�-�<˲�8]D�I[�E&��s/0��d�u8��er��PU5��� �B=V�.�Xu,H
��HS�=��Na*oǼx��D��������o�F�Fu�O8�Rվp;��m壉�Չ>XqL̪�x2]�I��̃��4�j 3�Y��͝F�Q��m�[��ɋC5Ts��AەN���+)��#�s�a��b�듵9^�p.b9Z��e�`�x}#]� ��!�HFd" �k��.��?���:�Ԓ�,�kܤT���ܐ���<��)i�:�S���K���3�*����j��j�B��B�^�@>f����V�߿��OD���|X$��]���i	yV�F��R����c{[��W#i���ʡ��t�zɑ�8�Fڐ��5��� �?�{�Ӧ������"������>};���9����,��bm� �Gf���
��<��S���^�s/����`n�43��="�2qc�d �\�A���)i���P�n������r��ř�o��i�!�fi�n�b��g1=^I��<��(zGͻ�La��+Ϯ��E��4ƌ�-n[��n����f�º�V�b���P쥫�L�\�fQ�3d��q��z�0Q��C����p��gi�bid0+�G��j�WH6��@稶��`�0\l�t����Upi7ƹܠ����_g$�ebmd�3��^��J�@��݌��N��r==��FqF���#gow���#L�5��߸0�h���%����-���dr���p!R�����v'��0�Z5=��j�oR�X5^0�����I�]�x�ʰ�tԦ�~��w����7�ȥ���"
��J� �Nn�KT	`����n��x��+����1�V�ʯ��`Z�&>�î�1��?5Ӳ�Y;�V`�/"���q���zp�`�3�벑���B��ܹ������\���7s����C(�`˧,��y��ڀi{5��a��`�	-�X���f� �	�O2D��Ѐ��֑��o� ��j&��4�0[9��t��
�%w]T��6��V֨��g���g��̈́��/�((��j��*��g^��>m�%���Q�3l��w��9�ǧ3����\hd	�{��6��g4G�,�0���Q�F��D��g*�ps��#=N1V!8ƭַ(]`QizP�G|z%?#&>v��nX ���쳀,5���[3	�F$����6p��*r��C���r@\����N��+͎���t�ʯNS
�Ƶ F�]� r �ƶ�̮]$֬�� �t1�=[���-�@IW���^x�M�&ԭ9�����rx�0r�%m&��o_�w���X�səm~��Zm�����I%�;�̓�'^�Oj��]=H��w��9�,oN0�;*;��"dܧ/`R7�����d��T� 1�pX�>��[�Pheg.APh]x��_kׅ������E�^�f\o���jY��	�S�5�!�N��4%GD�V��܇�����t��Yo��+����!�BrB�����_�S!W���'
�Z���4�,ǌK������M����#�0��5v����]�;1Y� �3�2~�G�&�m�δf��e�
W���(�<_��nj+$V|ztGu�&���1s�rw�b���$Im,}�\��VX�Eŀ�`Z���Q���5�-��CI�O">&z�$�0k���M��1*��N?����GZ^�"��g��*ն���ذ� �t��{ X38~MzW:m���A@d�G(�L֠7�qxT��5�={����T��G2ۗ� �ی��y9�'mp�[$f�n��[���PB�r#��E��m||eo���C���H!�АL%�E��{�hgog�yܱ��0������X���\���K-��|��}d�����C��O0��>�����^���&�tnl|y��s�	r�'��ûl���?̮��5D��ǰ�o]刟�'.���K�"��P��G'!���RF�	������a®x�l��Z�v��q ��pڒ��5bꪗ�{TX�`f�>=�,/�TU�Z:�O� ���y?�bP=��a�-�B�S���UuС� �"��`���B���W�%���k�i����DOK�f��`����d�wqo���\h�I�qQ���d�l���q�;���|U��¨��S�����]s���&Q�>qXp�4J5N��x*Y_%4wg_Pa���#��K�b�`�)}���JR���R&��r��ɢ�r�i"*"+|���ܡ#򪥑�4�Q1C���
���pZ�S�H�I#��?�X�j_4[V��U��i�����������u��I��z5-)����-CL�Γ�3��3�Yئ������f�%F5B]XjvL�ٛ��c��{m���d�������4*U�����	�
�)n�k�KyWBF� ;n��������Ȉ��!�n�ʕ�`�+��V���IX��I)U3 ?Ʀ���� �A��Ѕf==��^ݶQ��vu�ĻQ�}�fYH��)}�b,/�>��G��
���Ƴ��#b~�K �- ��@~���j�l�ڪ�*��"ʁ��y���'Ƌ ��q�3K)��l��[�����
�g��b���@�1W�62��;�9��z�r�t��ۆV+�"5������~#�$Ҏ�p���>f��(dM��ǿQ��r��vK0��yn� f�0@�r)F����o�^$��H�BT��B8����c�&�hU�ґ���T���' k&��o�mK�ܬv�v�@I35��v�e'��E?*�^�*�ێ�Nr����do���آ��Lr[fن8L���N8�v�{�q�2���y}̶rʆ��;s��~v�P�%aH��P~0Uc�6?�@�3Ι���K�*d�޺�$_+������� ��hᬑE���Z<�	onhDy�u+}%tI��!Ktw\�=Ȕ�t�ܯ��r�k�7�Z6K��oÐ�7��A`�T��%�7$z�"R+�Y�I%[�����6���gSECA�X��;7V�����z�=�N�6sK�{��R^(@k�T-�Ą��)���chVo;<D֛+��.[�M^6�_z9�.L^�+M�M���Bg�G�WԴORx�>\h̙�;q��X��k^����
����~�����4���d�a��6m�Z RlY�8�?!t᜙&���(�`*���WBA��ʍ��Q4mms�� ɇ�Q������^+�~\�{��V����n�;6ў�K�Զ||[^�?����yw�J?���(�,��,���:�>92��U��k��r�S:�X����#�{z(�k5Q�s!N⻺?������:!�^6��g�E��c����7��R2�{w�f{-?�׻����p�����Y2�XF���ӭ�e���ˆ|�I:E)+�[h��"�!�����l�$�!Zx�,J-܄u������	;8�vF��*g�Odr�q�:pH{0Q
/�Z#����[��5��lte���]ޔ��Z(׿�&�ܚN�Ä{g��B����y�tu�?���e��H��?��u7�B_�Q��8�q����:�,M��k�%{��Q�� _5�F%�n<N��@��|7�p:�q��i��\?���U�I ���Kw��EFv 90=C���G��d�w�!�E�.���eF��Us>���k��ǭO�jX��Z`W	��T���[c��?h��]U.�����V��(�K��[H�[�c�X�/<�н�R5��+�w�X�6:Q>%��mK���$#�e��_��߯D_Hd��w���٭ �r��h�
�X �f����7��}��	�_�2 L��}7����tsm�WGomfNR��W��"+X8�'���}�)�������H�~�7p���=���6�`�@m����X��h���1�.|7�P�B�C������X���M��� �{�K �[[Ԍ��e�n>� ����0T����E
 $0a��t�&Q2:	<O����L��d-$�[X�Іo��mX��'�#�
���lo2�S��N����E�-�FQ��UzIi|%�����@�	���O�.��Q��U{ā���Nꊎ�����V�v�HÔ؈�q7��&�+Xɕw�� @��y
�h(̃L!@���Kd��H��Z���a}�x�UÁ���������]@��F$�}Q��Y bP%P���GQ<wۈ/yt�0AH�%����N�qn$�fT��T������RY����WB���44b�����٪`.l��%��߿uД˜�ߟNV����S�1Lt�N��q��+	]��we�v�H��.�V��81�5��@
�w.l�����;�27S8aZ���S�(W����(Ln��� ��N������p|`y_`+�'���Y^��#| ����~	V�+����+8�6����h	>!�D����¢���9���:��킷b#�2ZǼ�C ~\t�-%-,�FM��1����9ġ#}��Y�l~w�9��PUk��]�R\�>����2�c!9�S�y���@~�CZ�Y�R
�@B-��H�gl���r��RPM��"+�4�3���;��j��5�7LT�L�